magic
tech sky130A
magscale 1 2
timestamp 1656859285
<< viali >>
rect 14565 69445 14599 69479
rect 19717 69445 19751 69479
rect 20821 69445 20855 69479
rect 35633 69445 35667 69479
rect 67649 69445 67683 69479
rect 1409 69377 1443 69411
rect 7849 69377 7883 69411
rect 46581 69377 46615 69411
rect 55505 69377 55539 69411
rect 57897 69377 57931 69411
rect 1593 69309 1627 69343
rect 65809 69309 65843 69343
rect 65993 69309 66027 69343
rect 14749 69241 14783 69275
rect 19901 69241 19935 69275
rect 21005 69241 21039 69275
rect 35909 69241 35943 69275
rect 2513 69173 2547 69207
rect 4813 69173 4847 69207
rect 6561 69173 6595 69207
rect 8033 69173 8067 69207
rect 11713 69173 11747 69207
rect 16865 69173 16899 69207
rect 24869 69173 24903 69207
rect 27353 69173 27387 69207
rect 31217 69173 31251 69207
rect 36645 69173 36679 69207
rect 37565 69173 37599 69207
rect 39037 69173 39071 69207
rect 41429 69173 41463 69207
rect 42901 69173 42935 69207
rect 45477 69173 45511 69207
rect 46121 69173 46155 69207
rect 46673 69173 46707 69207
rect 50721 69173 50755 69207
rect 52929 69173 52963 69207
rect 55689 69173 55723 69207
rect 56517 69173 56551 69207
rect 57345 69173 57379 69207
rect 57989 69173 58023 69207
rect 60657 69173 60691 69207
rect 62221 69173 62255 69207
rect 64429 69173 64463 69207
rect 65073 69173 65107 69207
rect 1409 68833 1443 68867
rect 2789 68833 2823 68867
rect 6009 68833 6043 68867
rect 6469 68833 6503 68867
rect 11069 68833 11103 68867
rect 11805 68833 11839 68867
rect 16129 68833 16163 68867
rect 16957 68833 16991 68867
rect 24685 68833 24719 68867
rect 25145 68833 25179 68867
rect 27077 68833 27111 68867
rect 27721 68833 27755 68867
rect 31033 68833 31067 68867
rect 31769 68833 31803 68867
rect 36277 68833 36311 68867
rect 36737 68833 36771 68867
rect 40325 68833 40359 68867
rect 41889 68833 41923 68867
rect 42625 68833 42659 68867
rect 43177 68833 43211 68867
rect 46397 68833 46431 68867
rect 46581 68833 46615 68867
rect 47041 68833 47075 68867
rect 50445 68833 50479 68867
rect 51549 68833 51583 68867
rect 52745 68833 52779 68867
rect 53205 68833 53239 68867
rect 56241 68833 56275 68867
rect 56701 68833 56735 68867
rect 60473 68833 60507 68867
rect 60933 68833 60967 68867
rect 62773 68833 62807 68867
rect 63233 68833 63267 68867
rect 66269 68833 66303 68867
rect 68109 68833 68143 68867
rect 4629 68765 4663 68799
rect 5365 68765 5399 68799
rect 10425 68765 10459 68799
rect 15485 68765 15519 68799
rect 38945 68765 38979 68799
rect 45293 68765 45327 68799
rect 48973 68765 49007 68799
rect 49433 68765 49467 68799
rect 59737 68765 59771 68799
rect 65625 68765 65659 68799
rect 1593 68697 1627 68731
rect 5457 68697 5491 68731
rect 6193 68697 6227 68731
rect 10517 68697 10551 68731
rect 11253 68697 11287 68731
rect 15577 68697 15611 68731
rect 16313 68697 16347 68731
rect 24869 68697 24903 68731
rect 27261 68697 27295 68731
rect 31217 68697 31251 68731
rect 36461 68697 36495 68731
rect 40509 68697 40543 68731
rect 42809 68697 42843 68731
rect 49525 68697 49559 68731
rect 50629 68697 50663 68731
rect 52929 68697 52963 68731
rect 56425 68697 56459 68731
rect 59829 68697 59863 68731
rect 60657 68697 60691 68731
rect 62957 68697 62991 68731
rect 66453 68697 66487 68731
rect 4721 68629 4755 68663
rect 39037 68629 39071 68663
rect 45385 68629 45419 68663
rect 65717 68629 65751 68663
rect 1869 68425 1903 68459
rect 24777 68425 24811 68459
rect 27261 68425 27295 68459
rect 31125 68425 31159 68459
rect 36553 68425 36587 68459
rect 42809 68425 42843 68459
rect 52837 68425 52871 68459
rect 56333 68425 56367 68459
rect 61669 68425 61703 68459
rect 39773 68357 39807 68391
rect 45385 68357 45419 68391
rect 58081 68357 58115 68391
rect 65717 68357 65751 68391
rect 1777 68289 1811 68323
rect 2513 68289 2547 68323
rect 24685 68289 24719 68323
rect 27169 68289 27203 68323
rect 31033 68289 31067 68323
rect 36461 68289 36495 68323
rect 37289 68289 37323 68323
rect 39589 68289 39623 68323
rect 42717 68289 42751 68323
rect 45201 68289 45235 68323
rect 49617 68289 49651 68323
rect 52745 68289 52779 68323
rect 56241 68289 56275 68323
rect 57897 68289 57931 68323
rect 61577 68289 61611 68323
rect 65533 68289 65567 68323
rect 3341 68221 3375 68255
rect 37473 68221 37507 68255
rect 38025 68221 38059 68255
rect 40049 68221 40083 68255
rect 45753 68221 45787 68255
rect 49801 68221 49835 68255
rect 50353 68221 50387 68255
rect 58357 68221 58391 68255
rect 65073 68221 65107 68255
rect 67005 68221 67039 68255
rect 37565 67881 37599 67915
rect 41429 67881 41463 67915
rect 50261 67881 50295 67915
rect 66269 67881 66303 67915
rect 67097 67881 67131 67915
rect 2329 67745 2363 67779
rect 4537 67745 4571 67779
rect 4721 67745 4755 67779
rect 5181 67745 5215 67779
rect 2053 67677 2087 67711
rect 37473 67677 37507 67711
rect 41337 67677 41371 67711
rect 50169 67677 50203 67711
rect 66177 67677 66211 67711
rect 67005 67677 67039 67711
rect 67741 67677 67775 67711
rect 68109 67609 68143 67643
rect 67649 67269 67683 67303
rect 1593 67201 1627 67235
rect 1869 67201 1903 67235
rect 2697 67201 2731 67235
rect 4353 67201 4387 67235
rect 3065 67133 3099 67167
rect 5181 67133 5215 67167
rect 65809 67133 65843 67167
rect 65993 67133 66027 67167
rect 67005 66793 67039 66827
rect 67557 66793 67591 66827
rect 2789 66657 2823 66691
rect 6009 66657 6043 66691
rect 1409 66589 1443 66623
rect 3985 66589 4019 66623
rect 5641 66589 5675 66623
rect 67465 66589 67499 66623
rect 1593 66521 1627 66555
rect 4997 66521 5031 66555
rect 1961 66249 1995 66283
rect 1869 66113 1903 66147
rect 2605 66113 2639 66147
rect 4353 66113 4387 66147
rect 36093 66113 36127 66147
rect 3709 66045 3743 66079
rect 5549 66045 5583 66079
rect 36369 66045 36403 66079
rect 65809 66045 65843 66079
rect 65993 66045 66027 66079
rect 67557 66045 67591 66079
rect 35909 65909 35943 65943
rect 36277 65909 36311 65943
rect 67005 65705 67039 65739
rect 67557 65705 67591 65739
rect 1685 65501 1719 65535
rect 2145 65501 2179 65535
rect 3249 65501 3283 65535
rect 3985 65501 4019 65535
rect 35173 65501 35207 65535
rect 35440 65501 35474 65535
rect 67465 65501 67499 65535
rect 2881 65433 2915 65467
rect 4813 65433 4847 65467
rect 2237 65365 2271 65399
rect 36553 65365 36587 65399
rect 1961 65093 1995 65127
rect 1777 65025 1811 65059
rect 4077 65025 4111 65059
rect 36093 65025 36127 65059
rect 36277 65025 36311 65059
rect 36369 65025 36403 65059
rect 38301 65025 38335 65059
rect 3617 64957 3651 64991
rect 4353 64957 4387 64991
rect 35909 64957 35943 64991
rect 38117 64821 38151 64855
rect 1961 64617 1995 64651
rect 37289 64617 37323 64651
rect 37473 64617 37507 64651
rect 36921 64549 36955 64583
rect 36277 64413 36311 64447
rect 37933 64413 37967 64447
rect 38200 64413 38234 64447
rect 36461 64345 36495 64379
rect 37289 64277 37323 64311
rect 39313 64277 39347 64311
rect 36737 64073 36771 64107
rect 37565 64073 37599 64107
rect 37933 64073 37967 64107
rect 36369 64005 36403 64039
rect 36585 64005 36619 64039
rect 34244 63937 34278 63971
rect 37749 63937 37783 63971
rect 38025 63937 38059 63971
rect 33977 63869 34011 63903
rect 35357 63733 35391 63767
rect 36553 63733 36587 63767
rect 67649 63733 67683 63767
rect 34713 63529 34747 63563
rect 36001 63529 36035 63563
rect 36737 63529 36771 63563
rect 37013 63393 37047 63427
rect 66269 63393 66303 63427
rect 1409 63325 1443 63359
rect 24501 63325 24535 63359
rect 34897 63325 34931 63359
rect 35633 63325 35667 63359
rect 36921 63325 36955 63359
rect 37105 63325 37139 63359
rect 37197 63325 37231 63359
rect 68109 63325 68143 63359
rect 1685 63257 1719 63291
rect 24869 63257 24903 63291
rect 66453 63257 66487 63291
rect 36001 63189 36035 63223
rect 36185 63189 36219 63223
rect 67557 62985 67591 63019
rect 28549 62917 28583 62951
rect 29285 62917 29319 62951
rect 35357 62917 35391 62951
rect 35557 62917 35591 62951
rect 23121 62849 23155 62883
rect 23489 62849 23523 62883
rect 24133 62849 24167 62883
rect 28457 62849 28491 62883
rect 34805 62849 34839 62883
rect 36185 62849 36219 62883
rect 36461 62849 36495 62883
rect 37657 62849 37691 62883
rect 37841 62849 37875 62883
rect 38557 62849 38591 62883
rect 67465 62849 67499 62883
rect 24501 62781 24535 62815
rect 29101 62781 29135 62815
rect 29561 62781 29595 62815
rect 32965 62781 32999 62815
rect 33149 62781 33183 62815
rect 36277 62781 36311 62815
rect 38301 62781 38335 62815
rect 35725 62713 35759 62747
rect 36645 62713 36679 62747
rect 35541 62645 35575 62679
rect 36185 62645 36219 62679
rect 37749 62645 37783 62679
rect 39681 62645 39715 62679
rect 33149 62441 33183 62475
rect 37749 62441 37783 62475
rect 23121 62305 23155 62339
rect 30849 62305 30883 62339
rect 35541 62305 35575 62339
rect 19901 62237 19935 62271
rect 22661 62237 22695 62271
rect 24409 62237 24443 62271
rect 26249 62237 26283 62271
rect 28089 62237 28123 62271
rect 29009 62237 29043 62271
rect 29745 62237 29779 62271
rect 30389 62237 30423 62271
rect 33057 62237 33091 62271
rect 35265 62237 35299 62271
rect 35357 62237 35391 62271
rect 38025 62237 38059 62271
rect 38117 62237 38151 62271
rect 38209 62237 38243 62271
rect 38393 62237 38427 62271
rect 67925 62237 67959 62271
rect 25329 62169 25363 62203
rect 26516 62169 26550 62203
rect 29837 62169 29871 62203
rect 30573 62169 30607 62203
rect 19901 62101 19935 62135
rect 27629 62101 27663 62135
rect 28273 62101 28307 62135
rect 28825 62101 28859 62135
rect 35541 62101 35575 62135
rect 26157 61897 26191 61931
rect 25145 61829 25179 61863
rect 27804 61829 27838 61863
rect 67649 61829 67683 61863
rect 19257 61761 19291 61795
rect 19513 61761 19547 61795
rect 21281 61761 21315 61795
rect 21833 61761 21867 61795
rect 25973 61761 26007 61795
rect 27537 61761 27571 61795
rect 29653 61761 29687 61795
rect 29920 61761 29954 61795
rect 33692 61761 33726 61795
rect 36001 61761 36035 61795
rect 36277 61761 36311 61795
rect 65809 61761 65843 61795
rect 22753 61693 22787 61727
rect 22937 61693 22971 61727
rect 23673 61693 23707 61727
rect 33425 61693 33459 61727
rect 35817 61693 35851 61727
rect 36093 61693 36127 61727
rect 36185 61693 36219 61727
rect 65993 61693 66027 61727
rect 20637 61557 20671 61591
rect 21097 61557 21131 61591
rect 21833 61557 21867 61591
rect 25237 61557 25271 61591
rect 28917 61557 28951 61591
rect 31033 61557 31067 61591
rect 34805 61557 34839 61591
rect 20729 61353 20763 61387
rect 23581 61353 23615 61387
rect 26433 61353 26467 61387
rect 28641 61353 28675 61387
rect 33057 61353 33091 61387
rect 67649 61353 67683 61387
rect 34805 61285 34839 61319
rect 19441 61217 19475 61251
rect 20361 61217 20395 61251
rect 21189 61217 21223 61251
rect 27721 61217 27755 61251
rect 19625 61149 19659 61183
rect 20545 61149 20579 61183
rect 21445 61149 21479 61183
rect 23489 61149 23523 61183
rect 24409 61149 24443 61183
rect 26617 61149 26651 61183
rect 27445 61149 27479 61183
rect 27537 61149 27571 61183
rect 28273 61149 28307 61183
rect 28457 61149 28491 61183
rect 30829 61149 30863 61183
rect 30922 61149 30956 61183
rect 31033 61149 31067 61183
rect 31217 61149 31251 61183
rect 31677 61149 31711 61183
rect 34989 61149 35023 61183
rect 35081 61149 35115 61183
rect 36001 61149 36035 61183
rect 36093 61149 36127 61183
rect 36185 61149 36219 61183
rect 36369 61149 36403 61183
rect 36829 61149 36863 61183
rect 38945 61149 38979 61183
rect 39865 61149 39899 61183
rect 67557 61149 67591 61183
rect 25237 61081 25271 61115
rect 30573 61081 30607 61115
rect 31922 61081 31956 61115
rect 34805 61081 34839 61115
rect 37074 61081 37108 61115
rect 38761 61081 38795 61115
rect 40132 61081 40166 61115
rect 19809 61013 19843 61047
rect 22569 61013 22603 61047
rect 35725 61013 35759 61047
rect 38209 61013 38243 61047
rect 41245 61013 41279 61047
rect 19533 60809 19567 60843
rect 26249 60809 26283 60843
rect 30297 60809 30331 60843
rect 36645 60809 36679 60843
rect 40049 60809 40083 60843
rect 1869 60741 1903 60775
rect 16129 60673 16163 60707
rect 17673 60673 17707 60707
rect 19717 60673 19751 60707
rect 22385 60673 22419 60707
rect 23489 60673 23523 60707
rect 25145 60673 25179 60707
rect 26433 60673 26467 60707
rect 27445 60673 27479 60707
rect 30573 60673 30607 60707
rect 30665 60673 30699 60707
rect 30778 60673 30812 60707
rect 30941 60673 30975 60707
rect 33701 60673 33735 60707
rect 35909 60673 35943 60707
rect 36553 60673 36587 60707
rect 36737 60673 36771 60707
rect 38117 60673 38151 60707
rect 38384 60673 38418 60707
rect 39957 60673 39991 60707
rect 40141 60673 40175 60707
rect 17417 60605 17451 60639
rect 22201 60605 22235 60639
rect 27261 60605 27295 60639
rect 27629 60605 27663 60639
rect 35725 60605 35759 60639
rect 65809 60605 65843 60639
rect 65993 60605 66027 60639
rect 67557 60605 67591 60639
rect 36093 60537 36127 60571
rect 2145 60469 2179 60503
rect 15945 60469 15979 60503
rect 18797 60469 18831 60503
rect 22569 60469 22603 60503
rect 23581 60469 23615 60503
rect 24961 60469 24995 60503
rect 33793 60469 33827 60503
rect 39497 60469 39531 60503
rect 25789 60265 25823 60299
rect 30389 60265 30423 60299
rect 31309 60265 31343 60299
rect 38761 60265 38795 60299
rect 39865 60265 39899 60299
rect 67373 60265 67407 60299
rect 68109 60265 68143 60299
rect 21465 60197 21499 60231
rect 17417 60129 17451 60163
rect 20821 60129 20855 60163
rect 21858 60129 21892 60163
rect 22017 60129 22051 60163
rect 27169 60129 27203 60163
rect 27813 60129 27847 60163
rect 28227 60129 28261 60163
rect 39129 60129 39163 60163
rect 42901 60129 42935 60163
rect 1869 60061 1903 60095
rect 15577 60061 15611 60095
rect 15844 60061 15878 60095
rect 17601 60061 17635 60095
rect 21005 60061 21039 60095
rect 21741 60061 21775 60095
rect 23765 60061 23799 60095
rect 23857 60061 23891 60095
rect 24409 60061 24443 60095
rect 24676 60061 24710 60095
rect 26341 60061 26375 60095
rect 27353 60061 27387 60095
rect 28089 60061 28123 60095
rect 28365 60061 28399 60095
rect 29745 60061 29779 60095
rect 30573 60061 30607 60095
rect 30849 60061 30883 60095
rect 31493 60061 31527 60095
rect 31769 60061 31803 60095
rect 32689 60061 32723 60095
rect 35541 60061 35575 60095
rect 38945 60061 38979 60095
rect 39221 60061 39255 60095
rect 40049 60061 40083 60095
rect 40141 60061 40175 60095
rect 67281 60061 67315 60095
rect 29009 59993 29043 60027
rect 32934 59993 32968 60027
rect 39865 59993 39899 60027
rect 43168 59993 43202 60027
rect 16957 59925 16991 59959
rect 17785 59925 17819 59959
rect 22661 59925 22695 59959
rect 26433 59925 26467 59959
rect 29561 59925 29595 59959
rect 30757 59925 30791 59959
rect 31677 59925 31711 59959
rect 34069 59925 34103 59959
rect 35357 59925 35391 59959
rect 44281 59925 44315 59959
rect 15853 59721 15887 59755
rect 17049 59721 17083 59755
rect 17693 59721 17727 59755
rect 22201 59721 22235 59755
rect 25513 59721 25547 59755
rect 28365 59721 28399 59755
rect 32229 59721 32263 59755
rect 36553 59721 36587 59755
rect 44097 59721 44131 59755
rect 23090 59653 23124 59687
rect 27230 59653 27264 59687
rect 33977 59653 34011 59687
rect 35633 59653 35667 59687
rect 1685 59585 1719 59619
rect 14657 59585 14691 59619
rect 15853 59585 15887 59619
rect 16865 59585 16899 59619
rect 17693 59585 17727 59619
rect 18613 59585 18647 59619
rect 18797 59585 18831 59619
rect 19533 59585 19567 59619
rect 22385 59585 22419 59619
rect 22845 59585 22879 59619
rect 25237 59585 25271 59619
rect 25329 59585 25363 59619
rect 26985 59585 27019 59619
rect 29644 59585 29678 59619
rect 32505 59585 32539 59619
rect 32597 59585 32631 59619
rect 32689 59585 32723 59619
rect 32873 59585 32907 59619
rect 33793 59585 33827 59619
rect 37545 59585 37579 59619
rect 39681 59585 39715 59619
rect 41429 59585 41463 59619
rect 41613 59585 41647 59619
rect 41705 59585 41739 59619
rect 43361 59585 43395 59619
rect 44005 59585 44039 59619
rect 44189 59585 44223 59619
rect 67281 59585 67315 59619
rect 1869 59517 1903 59551
rect 2789 59517 2823 59551
rect 16681 59517 16715 59551
rect 19650 59517 19684 59551
rect 19809 59517 19843 59551
rect 29377 59517 29411 59551
rect 36093 59517 36127 59551
rect 37289 59517 37323 59551
rect 39405 59517 39439 59551
rect 43177 59517 43211 59551
rect 43269 59517 43303 59551
rect 43453 59517 43487 59551
rect 19257 59449 19291 59483
rect 20453 59449 20487 59483
rect 36369 59449 36403 59483
rect 14473 59381 14507 59415
rect 24225 59381 24259 59415
rect 30757 59381 30791 59415
rect 38669 59381 38703 59415
rect 41429 59381 41463 59415
rect 42993 59381 43027 59415
rect 67373 59381 67407 59415
rect 2053 59177 2087 59211
rect 17417 59177 17451 59211
rect 29745 59177 29779 59211
rect 29929 59177 29963 59211
rect 31493 59177 31527 59211
rect 36277 59177 36311 59211
rect 39865 59177 39899 59211
rect 42257 59177 42291 59211
rect 42993 59177 43027 59211
rect 15485 59109 15519 59143
rect 38669 59041 38703 59075
rect 38945 59041 38979 59075
rect 39129 59041 39163 59075
rect 40141 59041 40175 59075
rect 40233 59041 40267 59075
rect 1961 58973 1995 59007
rect 14105 58973 14139 59007
rect 14372 58973 14406 59007
rect 17601 58973 17635 59007
rect 19441 58973 19475 59007
rect 20177 58973 20211 59007
rect 21649 58973 21683 59007
rect 25421 58973 25455 59007
rect 31677 58973 31711 59007
rect 31953 58973 31987 59007
rect 34897 58973 34931 59007
rect 37197 58973 37231 59007
rect 37381 58973 37415 59007
rect 38853 58973 38887 59007
rect 39037 58973 39071 59007
rect 40049 58973 40083 59007
rect 40325 58973 40359 59007
rect 40877 58973 40911 59007
rect 43177 58973 43211 59007
rect 43269 58973 43303 59007
rect 29561 58905 29595 58939
rect 35164 58905 35198 58939
rect 41144 58905 41178 58939
rect 42993 58905 43027 58939
rect 19441 58837 19475 58871
rect 19993 58837 20027 58871
rect 21465 58837 21499 58871
rect 25237 58837 25271 58871
rect 29771 58837 29805 58871
rect 31861 58837 31895 58871
rect 37565 58837 37599 58871
rect 14105 58633 14139 58667
rect 15117 58633 15151 58667
rect 20453 58633 20487 58667
rect 21113 58633 21147 58667
rect 21281 58633 21315 58667
rect 23213 58633 23247 58667
rect 25605 58633 25639 58667
rect 32505 58633 32539 58667
rect 37289 58633 37323 58667
rect 39957 58633 39991 58667
rect 41245 58633 41279 58667
rect 43269 58633 43303 58667
rect 19340 58565 19374 58599
rect 20913 58565 20947 58599
rect 22078 58565 22112 58599
rect 29745 58565 29779 58599
rect 38117 58565 38151 58599
rect 38301 58565 38335 58599
rect 39773 58565 39807 58599
rect 13921 58497 13955 58531
rect 14841 58497 14875 58531
rect 14933 58497 14967 58531
rect 17141 58497 17175 58531
rect 19073 58497 19107 58531
rect 24317 58497 24351 58531
rect 25329 58497 25363 58531
rect 25421 58497 25455 58531
rect 26341 58497 26375 58531
rect 27353 58497 27387 58531
rect 27905 58497 27939 58531
rect 28942 58497 28976 58531
rect 29101 58497 29135 58531
rect 30205 58497 30239 58531
rect 31309 58497 31343 58531
rect 32321 58497 32355 58531
rect 32597 58497 32631 58531
rect 33609 58497 33643 58531
rect 37473 58497 37507 58531
rect 39037 58497 39071 58531
rect 39221 58497 39255 58531
rect 40049 58497 40083 58531
rect 40509 58497 40543 58531
rect 41429 58497 41463 58531
rect 41705 58497 41739 58531
rect 43637 58497 43671 58531
rect 44465 58497 44499 58531
rect 21833 58429 21867 58463
rect 28089 58429 28123 58463
rect 28549 58429 28583 58463
rect 28825 58429 28859 58463
rect 39313 58429 39347 58463
rect 43453 58429 43487 58463
rect 43545 58429 43579 58463
rect 43729 58429 43763 58463
rect 44281 58429 44315 58463
rect 39773 58361 39807 58395
rect 16957 58293 16991 58327
rect 21097 58293 21131 58327
rect 24409 58293 24443 58327
rect 26341 58293 26375 58327
rect 27169 58293 27203 58327
rect 30389 58293 30423 58327
rect 31125 58293 31159 58327
rect 32137 58293 32171 58327
rect 33701 58293 33735 58327
rect 38853 58293 38887 58327
rect 40693 58293 40727 58327
rect 41613 58293 41647 58327
rect 44649 58293 44683 58327
rect 67649 58293 67683 58327
rect 19993 58089 20027 58123
rect 20177 58089 20211 58123
rect 21005 58089 21039 58123
rect 28089 58089 28123 58123
rect 38577 58021 38611 58055
rect 24593 57953 24627 57987
rect 26157 57953 26191 57987
rect 26709 57953 26743 57987
rect 15853 57885 15887 57919
rect 16037 57885 16071 57919
rect 16497 57885 16531 57919
rect 16764 57885 16798 57919
rect 20821 57885 20855 57919
rect 22477 57885 22511 57919
rect 24409 57885 24443 57919
rect 26976 57885 27010 57919
rect 29653 57885 29687 57919
rect 30297 57885 30331 57919
rect 30564 57885 30598 57919
rect 32413 57885 32447 57919
rect 34713 57885 34747 57919
rect 36921 57885 36955 57919
rect 38577 57885 38611 57919
rect 38761 57885 38795 57919
rect 44281 57885 44315 57919
rect 45017 57885 45051 57919
rect 66269 57885 66303 57919
rect 68109 57885 68143 57919
rect 19809 57817 19843 57851
rect 22744 57817 22778 57851
rect 29745 57817 29779 57851
rect 32658 57817 32692 57851
rect 34958 57817 34992 57851
rect 45262 57817 45296 57851
rect 66453 57817 66487 57851
rect 17877 57749 17911 57783
rect 20009 57749 20043 57783
rect 23857 57749 23891 57783
rect 31677 57749 31711 57783
rect 33793 57749 33827 57783
rect 36093 57749 36127 57783
rect 36737 57749 36771 57783
rect 44097 57749 44131 57783
rect 46397 57749 46431 57783
rect 17417 57545 17451 57579
rect 30941 57545 30975 57579
rect 39681 57545 39715 57579
rect 67557 57545 67591 57579
rect 22753 57477 22787 57511
rect 25136 57477 25170 57511
rect 27813 57477 27847 57511
rect 29929 57477 29963 57511
rect 30145 57477 30179 57511
rect 32137 57477 32171 57511
rect 33885 57477 33919 57511
rect 37657 57477 37691 57511
rect 39589 57477 39623 57511
rect 14648 57409 14682 57443
rect 17141 57409 17175 57443
rect 17233 57409 17267 57443
rect 18337 57409 18371 57443
rect 19190 57409 19224 57443
rect 23029 57409 23063 57443
rect 23121 57409 23155 57443
rect 23213 57409 23247 57443
rect 23397 57409 23431 57443
rect 24317 57409 24351 57443
rect 27629 57409 27663 57443
rect 30849 57409 30883 57443
rect 32413 57409 32447 57443
rect 32505 57409 32539 57443
rect 32597 57409 32631 57443
rect 32781 57409 32815 57443
rect 33701 57409 33735 57443
rect 36093 57409 36127 57443
rect 36185 57409 36219 57443
rect 37473 57409 37507 57443
rect 38853 57409 38887 57443
rect 41337 57409 41371 57443
rect 42717 57409 42751 57443
rect 67465 57409 67499 57443
rect 14381 57341 14415 57375
rect 18153 57341 18187 57375
rect 19073 57341 19107 57375
rect 19349 57341 19383 57375
rect 24409 57341 24443 57375
rect 24869 57341 24903 57375
rect 27445 57341 27479 57375
rect 34529 57341 34563 57375
rect 37289 57341 37323 57375
rect 38761 57341 38795 57375
rect 38945 57341 38979 57375
rect 42809 57341 42843 57375
rect 42901 57341 42935 57375
rect 15761 57273 15795 57307
rect 18797 57273 18831 57307
rect 26249 57273 26283 57307
rect 30297 57273 30331 57307
rect 19993 57205 20027 57239
rect 30113 57205 30147 57239
rect 36369 57205 36403 57239
rect 38577 57205 38611 57239
rect 41153 57205 41187 57239
rect 42533 57205 42567 57239
rect 14381 57001 14415 57035
rect 21649 57001 21683 57035
rect 24961 57001 24995 57035
rect 28181 57001 28215 57035
rect 33977 57001 34011 57035
rect 37657 57001 37691 57035
rect 39129 57001 39163 57035
rect 44465 57001 44499 57035
rect 35357 56933 35391 56967
rect 15025 56865 15059 56899
rect 18429 56865 18463 56899
rect 36277 56865 36311 56899
rect 40785 56865 40819 56899
rect 43085 56865 43119 56899
rect 1409 56797 1443 56831
rect 14197 56797 14231 56831
rect 15209 56797 15243 56831
rect 17141 56797 17175 56831
rect 18153 56797 18187 56831
rect 18245 56797 18279 56831
rect 19625 56797 19659 56831
rect 20545 56797 20579 56831
rect 21833 56797 21867 56831
rect 22109 56797 22143 56831
rect 26157 56797 26191 56831
rect 30849 56797 30883 56831
rect 33517 56797 33551 56831
rect 34161 56797 34195 56831
rect 36544 56797 36578 56831
rect 38945 56797 38979 56831
rect 45385 56797 45419 56831
rect 46857 56797 46891 56831
rect 50353 56797 50387 56831
rect 67649 56797 67683 56831
rect 24869 56729 24903 56763
rect 26424 56729 26458 56763
rect 28089 56729 28123 56763
rect 31116 56729 31150 56763
rect 35173 56729 35207 56763
rect 38577 56729 38611 56763
rect 41052 56729 41086 56763
rect 43352 56729 43386 56763
rect 47124 56729 47158 56763
rect 67925 56729 67959 56763
rect 1593 56661 1627 56695
rect 15393 56661 15427 56695
rect 16957 56661 16991 56695
rect 19809 56661 19843 56695
rect 20361 56661 20395 56695
rect 22017 56661 22051 56695
rect 27537 56661 27571 56695
rect 32229 56661 32263 56695
rect 33333 56661 33367 56695
rect 38761 56661 38795 56695
rect 38853 56661 38887 56695
rect 42165 56661 42199 56695
rect 45385 56661 45419 56695
rect 48237 56661 48271 56695
rect 50169 56661 50203 56695
rect 67281 56661 67315 56695
rect 26157 56457 26191 56491
rect 30849 56457 30883 56491
rect 35817 56457 35851 56491
rect 40877 56457 40911 56491
rect 43361 56457 43395 56491
rect 16948 56389 16982 56423
rect 19984 56389 20018 56423
rect 33578 56389 33612 56423
rect 35449 56389 35483 56423
rect 49424 56389 49458 56423
rect 15117 56321 15151 56355
rect 19717 56321 19751 56355
rect 22017 56321 22051 56355
rect 22201 56321 22235 56355
rect 22293 56321 22327 56355
rect 24777 56321 24811 56355
rect 25513 56321 25547 56355
rect 26157 56321 26191 56355
rect 27436 56321 27470 56355
rect 35541 56321 35575 56355
rect 35633 56321 35667 56355
rect 36369 56321 36403 56355
rect 39221 56321 39255 56355
rect 39313 56321 39347 56355
rect 39405 56321 39439 56355
rect 40509 56321 40543 56355
rect 40693 56321 40727 56355
rect 42625 56321 42659 56355
rect 43545 56321 43579 56355
rect 45201 56321 45235 56355
rect 45468 56321 45502 56355
rect 48237 56321 48271 56355
rect 48329 56321 48363 56355
rect 16681 56253 16715 56287
rect 27169 56253 27203 56287
rect 29009 56253 29043 56287
rect 29193 56253 29227 56287
rect 29929 56253 29963 56287
rect 30067 56253 30101 56287
rect 30205 56253 30239 56287
rect 33333 56253 33367 56287
rect 42901 56253 42935 56287
rect 43821 56253 43855 56287
rect 49157 56253 49191 56287
rect 14933 56185 14967 56219
rect 18061 56185 18095 56219
rect 28549 56185 28583 56219
rect 29653 56185 29687 56219
rect 35265 56185 35299 56219
rect 39037 56185 39071 56219
rect 39589 56185 39623 56219
rect 43729 56185 43763 56219
rect 21097 56117 21131 56151
rect 21833 56117 21867 56151
rect 24593 56117 24627 56151
rect 25329 56117 25363 56151
rect 34713 56117 34747 56151
rect 36553 56117 36587 56151
rect 42441 56117 42475 56151
rect 42809 56117 42843 56151
rect 46581 56117 46615 56151
rect 48513 56117 48547 56151
rect 50537 56117 50571 56151
rect 16037 55913 16071 55947
rect 20085 55913 20119 55947
rect 20269 55913 20303 55947
rect 23213 55913 23247 55947
rect 26525 55913 26559 55947
rect 30573 55913 30607 55947
rect 31217 55913 31251 55947
rect 45845 55913 45879 55947
rect 46857 55913 46891 55947
rect 48789 55913 48823 55947
rect 50537 55913 50571 55947
rect 29929 55845 29963 55879
rect 36921 55845 36955 55879
rect 38209 55845 38243 55879
rect 24501 55777 24535 55811
rect 27537 55777 27571 55811
rect 28457 55777 28491 55811
rect 36461 55777 36495 55811
rect 38853 55777 38887 55811
rect 45017 55777 45051 55811
rect 47685 55777 47719 55811
rect 50169 55777 50203 55811
rect 14841 55709 14875 55743
rect 16037 55709 16071 55743
rect 16773 55709 16807 55743
rect 21833 55709 21867 55743
rect 24768 55709 24802 55743
rect 26709 55709 26743 55743
rect 27261 55709 27295 55743
rect 27353 55709 27387 55743
rect 28641 55709 28675 55743
rect 29745 55709 29779 55743
rect 31217 55709 31251 55743
rect 32321 55709 32355 55743
rect 36001 55709 36035 55743
rect 36369 55709 36403 55743
rect 37105 55709 37139 55743
rect 37473 55709 37507 55743
rect 38209 55709 38243 55743
rect 38945 55709 38979 55743
rect 39037 55709 39071 55743
rect 40141 55709 40175 55743
rect 45201 55709 45235 55743
rect 45385 55709 45419 55743
rect 46029 55709 46063 55743
rect 46857 55709 46891 55743
rect 47593 55709 47627 55743
rect 48605 55709 48639 55743
rect 50353 55709 50387 55743
rect 19901 55641 19935 55675
rect 22100 55641 22134 55675
rect 30389 55641 30423 55675
rect 32505 55641 32539 55675
rect 34161 55641 34195 55675
rect 37289 55641 37323 55675
rect 37933 55641 37967 55675
rect 38117 55641 38151 55675
rect 40408 55641 40442 55675
rect 47869 55641 47903 55675
rect 14657 55573 14691 55607
rect 16773 55573 16807 55607
rect 20101 55573 20135 55607
rect 25881 55573 25915 55607
rect 28825 55573 28859 55607
rect 30589 55573 30623 55607
rect 30757 55573 30791 55607
rect 35725 55573 35759 55607
rect 36093 55573 36127 55607
rect 36185 55573 36219 55607
rect 37197 55573 37231 55607
rect 38669 55573 38703 55607
rect 41521 55573 41555 55607
rect 47593 55573 47627 55607
rect 25421 55369 25455 55403
rect 27721 55369 27755 55403
rect 28549 55369 28583 55403
rect 31401 55369 31435 55403
rect 32689 55369 32723 55403
rect 36645 55369 36679 55403
rect 40509 55369 40543 55403
rect 43913 55369 43947 55403
rect 47593 55369 47627 55403
rect 14464 55301 14498 55335
rect 37749 55301 37783 55335
rect 13645 55233 13679 55267
rect 16957 55233 16991 55267
rect 17224 55233 17258 55267
rect 18981 55233 19015 55267
rect 23305 55233 23339 55267
rect 25145 55233 25179 55267
rect 25237 55233 25271 55267
rect 27629 55233 27663 55267
rect 28733 55233 28767 55267
rect 31585 55233 31619 55267
rect 32597 55233 32631 55267
rect 33609 55233 33643 55267
rect 33876 55233 33910 55267
rect 35817 55233 35851 55267
rect 36001 55233 36035 55267
rect 36553 55233 36587 55267
rect 38945 55233 38979 55267
rect 39129 55233 39163 55267
rect 40693 55233 40727 55267
rect 42533 55233 42567 55267
rect 42800 55233 42834 55267
rect 45845 55233 45879 55267
rect 47777 55233 47811 55267
rect 48513 55233 48547 55267
rect 50353 55233 50387 55267
rect 51273 55233 51307 55267
rect 13737 55165 13771 55199
rect 14197 55165 14231 55199
rect 18797 55165 18831 55199
rect 23581 55165 23615 55199
rect 39221 55165 39255 55199
rect 40969 55165 41003 55199
rect 38761 55097 38795 55131
rect 40877 55097 40911 55131
rect 15577 55029 15611 55063
rect 18337 55029 18371 55063
rect 19165 55029 19199 55063
rect 34989 55029 35023 55063
rect 35817 55029 35851 55063
rect 37841 55029 37875 55063
rect 45753 55029 45787 55063
rect 48329 55029 48363 55063
rect 50353 55029 50387 55063
rect 51089 55029 51123 55063
rect 15301 54825 15335 54859
rect 17693 54825 17727 54859
rect 21741 54825 21775 54859
rect 34713 54825 34747 54859
rect 35081 54825 35115 54859
rect 38669 54825 38703 54859
rect 45201 54825 45235 54859
rect 20821 54757 20855 54791
rect 31401 54757 31435 54791
rect 35633 54757 35667 54791
rect 32597 54689 32631 54723
rect 45753 54689 45787 54723
rect 50445 54689 50479 54723
rect 15025 54621 15059 54655
rect 15117 54621 15151 54655
rect 17877 54621 17911 54655
rect 19625 54621 19659 54655
rect 20361 54621 20395 54655
rect 21005 54621 21039 54655
rect 21281 54621 21315 54655
rect 22017 54621 22051 54655
rect 22109 54621 22143 54655
rect 22201 54621 22235 54655
rect 22385 54621 22419 54655
rect 23213 54621 23247 54655
rect 23305 54621 23339 54655
rect 23397 54621 23431 54655
rect 23581 54621 23615 54655
rect 25421 54621 25455 54655
rect 29009 54621 29043 54655
rect 30113 54621 30147 54655
rect 31585 54621 31619 54655
rect 31769 54621 31803 54655
rect 31861 54621 31895 54655
rect 34897 54621 34931 54655
rect 35173 54621 35207 54655
rect 35817 54621 35851 54655
rect 35909 54621 35943 54655
rect 38485 54621 38519 54655
rect 38761 54621 38795 54655
rect 42993 54621 43027 54655
rect 44189 54621 44223 54655
rect 45017 54621 45051 54655
rect 47685 54621 47719 54655
rect 47952 54621 47986 54655
rect 50712 54621 50746 54655
rect 21189 54553 21223 54587
rect 28825 54553 28859 54587
rect 32413 54553 32447 54587
rect 35633 54553 35667 54587
rect 43177 54553 43211 54587
rect 45998 54553 46032 54587
rect 19625 54485 19659 54519
rect 20177 54485 20211 54519
rect 22937 54485 22971 54519
rect 25237 54485 25271 54519
rect 30113 54485 30147 54519
rect 38301 54485 38335 54519
rect 44281 54485 44315 54519
rect 47133 54485 47167 54519
rect 49065 54485 49099 54519
rect 51825 54485 51859 54519
rect 33517 54281 33551 54315
rect 45661 54281 45695 54315
rect 47777 54281 47811 54315
rect 48973 54281 49007 54315
rect 50261 54281 50295 54315
rect 19165 54213 19199 54247
rect 19892 54213 19926 54247
rect 21833 54213 21867 54247
rect 22201 54213 22235 54247
rect 37832 54213 37866 54247
rect 6377 54145 6411 54179
rect 15945 54145 15979 54179
rect 17325 54145 17359 54179
rect 18245 54145 18279 54179
rect 19625 54145 19659 54179
rect 22017 54145 22051 54179
rect 22293 54145 22327 54179
rect 23213 54145 23247 54179
rect 23469 54145 23503 54179
rect 25053 54145 25087 54179
rect 26341 54145 26375 54179
rect 27241 54145 27275 54179
rect 29837 54145 29871 54179
rect 30104 54145 30138 54179
rect 32404 54145 32438 54179
rect 37565 54145 37599 54179
rect 40049 54145 40083 54179
rect 40141 54145 40175 54179
rect 40325 54145 40359 54179
rect 40969 54145 41003 54179
rect 41429 54145 41463 54179
rect 43637 54145 43671 54179
rect 43893 54145 43927 54179
rect 45845 54145 45879 54179
rect 47593 54145 47627 54179
rect 48697 54145 48731 54179
rect 48789 54145 48823 54179
rect 50077 54145 50111 54179
rect 50905 54145 50939 54179
rect 6561 54077 6595 54111
rect 6929 54077 6963 54111
rect 15761 54077 15795 54111
rect 17509 54077 17543 54111
rect 18362 54077 18396 54111
rect 18521 54077 18555 54111
rect 26433 54077 26467 54111
rect 26985 54077 27019 54111
rect 32137 54077 32171 54111
rect 46121 54077 46155 54111
rect 49893 54077 49927 54111
rect 17969 54009 18003 54043
rect 24593 54009 24627 54043
rect 1961 53941 1995 53975
rect 16129 53941 16163 53975
rect 21005 53941 21039 53975
rect 25053 53941 25087 53975
rect 28365 53941 28399 53975
rect 31217 53941 31251 53975
rect 38945 53941 38979 53975
rect 40785 53941 40819 53975
rect 41521 53941 41555 53975
rect 45017 53941 45051 53975
rect 46029 53941 46063 53975
rect 50721 53941 50755 53975
rect 6101 53737 6135 53771
rect 16957 53737 16991 53771
rect 19993 53737 20027 53771
rect 20177 53737 20211 53771
rect 21557 53737 21591 53771
rect 26985 53737 27019 53771
rect 30021 53737 30055 53771
rect 30665 53737 30699 53771
rect 32873 53737 32907 53771
rect 43637 53737 43671 53771
rect 45293 53737 45327 53771
rect 48697 53737 48731 53771
rect 26249 53669 26283 53703
rect 48605 53669 48639 53703
rect 1409 53601 1443 53635
rect 2789 53601 2823 53635
rect 22753 53601 22787 53635
rect 24869 53601 24903 53635
rect 27997 53601 28031 53635
rect 31585 53601 31619 53635
rect 31861 53601 31895 53635
rect 35081 53601 35115 53635
rect 41521 53601 41555 53635
rect 6009 53533 6043 53567
rect 13461 53533 13495 53567
rect 14565 53533 14599 53567
rect 14657 53533 14691 53567
rect 15577 53533 15611 53567
rect 17417 53533 17451 53567
rect 21741 53533 21775 53567
rect 22017 53533 22051 53567
rect 22477 53533 22511 53567
rect 25136 53533 25170 53567
rect 27169 53533 27203 53567
rect 27721 53533 27755 53567
rect 27813 53533 27847 53567
rect 30849 53533 30883 53567
rect 33149 53533 33183 53567
rect 33241 53533 33275 53567
rect 33333 53533 33367 53567
rect 33517 53533 33551 53567
rect 35265 53533 35299 53567
rect 35541 53533 35575 53567
rect 36553 53533 36587 53567
rect 39221 53533 39255 53567
rect 40693 53533 40727 53567
rect 43637 53533 43671 53567
rect 43821 53533 43855 53567
rect 45109 53533 45143 53567
rect 46213 53533 46247 53567
rect 46397 53533 46431 53567
rect 48513 53533 48547 53567
rect 48789 53533 48823 53567
rect 50537 53533 50571 53567
rect 50804 53533 50838 53567
rect 20039 53499 20073 53533
rect 30067 53499 30101 53533
rect 1593 53465 1627 53499
rect 15844 53465 15878 53499
rect 18521 53465 18555 53499
rect 19809 53465 19843 53499
rect 21925 53465 21959 53499
rect 29837 53465 29871 53499
rect 35449 53465 35483 53499
rect 36820 53465 36854 53499
rect 40325 53465 40359 53499
rect 41788 53465 41822 53499
rect 48329 53465 48363 53499
rect 13461 53397 13495 53431
rect 14841 53397 14875 53431
rect 17601 53397 17635 53431
rect 18613 53397 18647 53431
rect 30205 53397 30239 53431
rect 37933 53397 37967 53431
rect 39221 53397 39255 53431
rect 42901 53397 42935 53431
rect 46397 53397 46431 53431
rect 48881 53397 48915 53431
rect 51917 53397 51951 53431
rect 2421 53193 2455 53227
rect 15761 53193 15795 53227
rect 16681 53193 16715 53227
rect 25697 53193 25731 53227
rect 29929 53193 29963 53227
rect 34529 53193 34563 53227
rect 35725 53193 35759 53227
rect 37289 53193 37323 53227
rect 40877 53193 40911 53227
rect 41521 53193 41555 53227
rect 41797 53193 41831 53227
rect 43453 53193 43487 53227
rect 45569 53193 45603 53227
rect 50261 53193 50295 53227
rect 50905 53193 50939 53227
rect 35357 53125 35391 53159
rect 35817 53125 35851 53159
rect 39764 53125 39798 53159
rect 41429 53125 41463 53159
rect 42441 53125 42475 53159
rect 43361 53125 43395 53159
rect 46489 53125 46523 53159
rect 2329 53057 2363 53091
rect 13553 53057 13587 53091
rect 13820 53057 13854 53091
rect 15761 53057 15795 53091
rect 16865 53057 16899 53091
rect 19533 53057 19567 53091
rect 20821 53057 20855 53091
rect 22661 53057 22695 53091
rect 24409 53057 24443 53091
rect 25421 53057 25455 53091
rect 25513 53057 25547 53091
rect 27629 53057 27663 53091
rect 29126 53057 29160 53091
rect 31125 53057 31159 53091
rect 33416 53057 33450 53091
rect 35633 53057 35667 53091
rect 37473 53057 37507 53091
rect 37749 53057 37783 53091
rect 39497 53057 39531 53091
rect 41326 53057 41360 53091
rect 41797 53057 41831 53091
rect 42625 53057 42659 53091
rect 42717 53057 42751 53091
rect 45477 53057 45511 53091
rect 45661 53057 45695 53091
rect 46305 53057 46339 53091
rect 46581 53057 46615 53091
rect 47869 53057 47903 53091
rect 47958 53060 47992 53094
rect 48053 53063 48087 53097
rect 48237 53057 48271 53091
rect 49893 53057 49927 53091
rect 50077 53057 50111 53091
rect 50721 53057 50755 53091
rect 22385 52989 22419 53023
rect 24685 52989 24719 53023
rect 28089 52989 28123 53023
rect 28273 52989 28307 53023
rect 29009 52989 29043 53023
rect 29285 52989 29319 53023
rect 33149 52989 33183 53023
rect 36093 52989 36127 53023
rect 47593 52989 47627 53023
rect 21005 52921 21039 52955
rect 28733 52921 28767 52955
rect 37657 52921 37691 52955
rect 42441 52921 42475 52955
rect 1777 52853 1811 52887
rect 14933 52853 14967 52887
rect 19349 52853 19383 52887
rect 27445 52853 27479 52887
rect 30941 52853 30975 52887
rect 36001 52853 36035 52887
rect 41705 52853 41739 52887
rect 46121 52853 46155 52887
rect 14105 52649 14139 52683
rect 16129 52649 16163 52683
rect 28181 52649 28215 52683
rect 29009 52649 29043 52683
rect 29745 52649 29779 52683
rect 33609 52649 33643 52683
rect 35449 52649 35483 52683
rect 43729 52649 43763 52683
rect 46489 52649 46523 52683
rect 24685 52581 24719 52615
rect 30573 52581 30607 52615
rect 35081 52581 35115 52615
rect 35633 52581 35667 52615
rect 46673 52581 46707 52615
rect 1409 52513 1443 52547
rect 1869 52513 1903 52547
rect 16957 52513 16991 52547
rect 18337 52513 18371 52547
rect 19349 52513 19383 52547
rect 28641 52513 28675 52547
rect 44373 52513 44407 52547
rect 14289 52445 14323 52479
rect 16681 52445 16715 52479
rect 18061 52445 18095 52479
rect 18153 52445 18187 52479
rect 21649 52445 21683 52479
rect 21738 52445 21772 52479
rect 21838 52445 21872 52479
rect 22017 52445 22051 52479
rect 22477 52445 22511 52479
rect 24501 52445 24535 52479
rect 25421 52445 25455 52479
rect 26801 52445 26835 52479
rect 27068 52445 27102 52479
rect 28825 52445 28859 52479
rect 29561 52445 29595 52479
rect 30389 52445 30423 52479
rect 31125 52445 31159 52479
rect 31381 52445 31415 52479
rect 33793 52445 33827 52479
rect 46121 52445 46155 52479
rect 46489 52445 46523 52479
rect 47593 52445 47627 52479
rect 50169 52445 50203 52479
rect 1593 52377 1627 52411
rect 16037 52377 16071 52411
rect 19594 52377 19628 52411
rect 21373 52377 21407 52411
rect 22744 52377 22778 52411
rect 35449 52377 35483 52411
rect 45477 52377 45511 52411
rect 45661 52377 45695 52411
rect 20729 52309 20763 52343
rect 23857 52309 23891 52343
rect 25237 52309 25271 52343
rect 32505 52309 32539 52343
rect 44097 52309 44131 52343
rect 44189 52309 44223 52343
rect 47777 52309 47811 52343
rect 50353 52309 50387 52343
rect 2053 52105 2087 52139
rect 19717 52037 19751 52071
rect 19933 52037 19967 52071
rect 22078 52037 22112 52071
rect 23673 52037 23707 52071
rect 32137 52037 32171 52071
rect 35173 52037 35207 52071
rect 35389 52037 35423 52071
rect 41521 52037 41555 52071
rect 45845 52037 45879 52071
rect 47838 52037 47872 52071
rect 32367 52003 32401 52037
rect 1961 51969 1995 52003
rect 14648 51969 14682 52003
rect 18337 51969 18371 52003
rect 20821 51969 20855 52003
rect 23949 51969 23983 52003
rect 24041 51969 24075 52003
rect 24133 51969 24167 52003
rect 24317 51969 24351 52003
rect 25145 51969 25179 52003
rect 25421 51969 25455 52003
rect 28089 51969 28123 52003
rect 28181 51969 28215 52003
rect 29653 51969 29687 52003
rect 30941 51969 30975 52003
rect 37841 51969 37875 52003
rect 38097 51969 38131 52003
rect 41245 51969 41279 52003
rect 41613 51969 41647 52003
rect 42441 51969 42475 52003
rect 43729 51969 43763 52003
rect 46121 51969 46155 52003
rect 46213 51969 46247 52003
rect 46305 51969 46339 52003
rect 46489 51969 46523 52003
rect 47593 51969 47627 52003
rect 49801 51969 49835 52003
rect 50068 51969 50102 52003
rect 67189 51969 67223 52003
rect 14381 51901 14415 51935
rect 17417 51901 17451 51935
rect 17601 51901 17635 51935
rect 18454 51901 18488 51935
rect 18613 51901 18647 51935
rect 19257 51901 19291 51935
rect 21833 51901 21867 51935
rect 29377 51901 29411 51935
rect 30665 51901 30699 51935
rect 41730 51901 41764 51935
rect 43821 51901 43855 51935
rect 18061 51833 18095 51867
rect 21005 51833 21039 51867
rect 32505 51833 32539 51867
rect 35541 51833 35575 51867
rect 39221 51833 39255 51867
rect 41889 51833 41923 51867
rect 48973 51833 49007 51867
rect 15761 51765 15795 51799
rect 19901 51765 19935 51799
rect 20085 51765 20119 51799
rect 23213 51765 23247 51799
rect 28365 51765 28399 51799
rect 32321 51765 32355 51799
rect 35357 51765 35391 51799
rect 42533 51765 42567 51799
rect 42901 51765 42935 51799
rect 43913 51765 43947 51799
rect 44097 51765 44131 51799
rect 51181 51765 51215 51799
rect 67281 51765 67315 51799
rect 15025 51561 15059 51595
rect 18153 51561 18187 51595
rect 19717 51561 19751 51595
rect 26801 51561 26835 51595
rect 31401 51561 31435 51595
rect 37381 51561 37415 51595
rect 41245 51561 41279 51595
rect 26249 51493 26283 51527
rect 36001 51493 36035 51527
rect 36461 51493 36495 51527
rect 51089 51493 51123 51527
rect 16037 51425 16071 51459
rect 20729 51425 20763 51459
rect 21557 51425 21591 51459
rect 29561 51425 29595 51459
rect 30205 51425 30239 51459
rect 30598 51425 30632 51459
rect 30757 51425 30791 51459
rect 38485 51425 38519 51459
rect 42533 51425 42567 51459
rect 49065 51425 49099 51459
rect 50261 51425 50295 51459
rect 66269 51425 66303 51459
rect 14197 51357 14231 51391
rect 15209 51357 15243 51391
rect 15761 51357 15795 51391
rect 15853 51357 15887 51391
rect 16773 51357 16807 51391
rect 19901 51357 19935 51391
rect 21833 51357 21867 51391
rect 23765 51357 23799 51391
rect 23857 51357 23891 51391
rect 24869 51357 24903 51391
rect 25136 51357 25170 51391
rect 26709 51357 26743 51391
rect 27997 51357 28031 51391
rect 28273 51357 28307 51391
rect 29745 51357 29779 51391
rect 30481 51357 30515 51391
rect 32781 51357 32815 51391
rect 34713 51357 34747 51391
rect 34897 51357 34931 51391
rect 35725 51357 35759 51391
rect 35817 51357 35851 51391
rect 36461 51357 36495 51391
rect 36737 51357 36771 51391
rect 37657 51357 37691 51391
rect 37749 51357 37783 51391
rect 37841 51357 37875 51391
rect 38025 51357 38059 51391
rect 38669 51357 38703 51391
rect 38853 51357 38887 51391
rect 38945 51357 38979 51391
rect 39865 51357 39899 51391
rect 40132 51357 40166 51391
rect 42349 51357 42383 51391
rect 42625 51357 42659 51391
rect 42993 51357 43027 51391
rect 43729 51357 43763 51391
rect 43821 51357 43855 51391
rect 44005 51357 44039 51391
rect 44097 51357 44131 51391
rect 45017 51357 45051 51391
rect 45201 51357 45235 51391
rect 46029 51357 46063 51391
rect 46213 51357 46247 51391
rect 48789 51357 48823 51391
rect 50445 51357 50479 51391
rect 50629 51357 50663 51391
rect 51273 51357 51307 51391
rect 17040 51289 17074 51323
rect 20545 51289 20579 51323
rect 33048 51289 33082 51323
rect 34805 51289 34839 51323
rect 35449 51289 35483 51323
rect 42901 51289 42935 51323
rect 66453 51289 66487 51323
rect 68109 51289 68143 51323
rect 14381 51221 14415 51255
rect 34161 51221 34195 51255
rect 35633 51221 35667 51255
rect 36645 51221 36679 51255
rect 43545 51221 43579 51255
rect 45109 51221 45143 51255
rect 46121 51221 46155 51255
rect 14105 51017 14139 51051
rect 16865 51017 16899 51051
rect 17417 51017 17451 51051
rect 21097 51017 21131 51051
rect 23673 51017 23707 51051
rect 24593 51017 24627 51051
rect 25697 51017 25731 51051
rect 28365 51017 28399 51051
rect 46397 51017 46431 51051
rect 46489 51017 46523 51051
rect 66453 51017 66487 51051
rect 31125 50949 31159 50983
rect 34437 50949 34471 50983
rect 35541 50949 35575 50983
rect 35757 50949 35791 50983
rect 46121 50949 46155 50983
rect 46305 50949 46339 50983
rect 14013 50881 14047 50915
rect 14657 50881 14691 50915
rect 16865 50881 16899 50915
rect 17601 50881 17635 50915
rect 19717 50881 19751 50915
rect 21005 50881 21039 50915
rect 23581 50881 23615 50915
rect 24501 50881 24535 50915
rect 25421 50881 25455 50915
rect 25513 50881 25547 50915
rect 26249 50881 26283 50915
rect 27252 50881 27286 50915
rect 29837 50881 29871 50915
rect 29929 50881 29963 50915
rect 30849 50881 30883 50915
rect 34161 50881 34195 50915
rect 36461 50881 36495 50915
rect 37749 50881 37783 50915
rect 38577 50881 38611 50915
rect 39497 50881 39531 50915
rect 40500 50881 40534 50915
rect 43729 50881 43763 50915
rect 43913 50881 43947 50915
rect 45109 50881 45143 50915
rect 46673 50881 46707 50915
rect 47685 50881 47719 50915
rect 48513 50881 48547 50915
rect 49893 50881 49927 50915
rect 50169 50881 50203 50915
rect 51457 50881 51491 50915
rect 51641 50881 51675 50915
rect 52929 50881 52963 50915
rect 66361 50881 66395 50915
rect 26433 50813 26467 50847
rect 26985 50813 27019 50847
rect 34437 50813 34471 50847
rect 39773 50813 39807 50847
rect 40233 50813 40267 50847
rect 43821 50813 43855 50847
rect 44005 50813 44039 50847
rect 44833 50813 44867 50847
rect 48789 50813 48823 50847
rect 51273 50813 51307 50847
rect 34253 50745 34287 50779
rect 35909 50745 35943 50779
rect 36645 50745 36679 50779
rect 38025 50745 38059 50779
rect 38669 50745 38703 50779
rect 41613 50745 41647 50779
rect 43545 50745 43579 50779
rect 14749 50677 14783 50711
rect 19533 50677 19567 50711
rect 30113 50677 30147 50711
rect 35725 50677 35759 50711
rect 47593 50677 47627 50711
rect 48605 50677 48639 50711
rect 49065 50677 49099 50711
rect 52745 50677 52779 50711
rect 27629 50473 27663 50507
rect 32505 50473 32539 50507
rect 41061 50473 41095 50507
rect 41429 50473 41463 50507
rect 47317 50473 47351 50507
rect 50353 50473 50387 50507
rect 52929 50473 52963 50507
rect 45661 50405 45695 50439
rect 50721 50405 50755 50439
rect 21097 50337 21131 50371
rect 24409 50337 24443 50371
rect 41521 50337 41555 50371
rect 47133 50337 47167 50371
rect 12633 50269 12667 50303
rect 15117 50269 15151 50303
rect 15209 50269 15243 50303
rect 17049 50269 17083 50303
rect 19257 50269 19291 50303
rect 19524 50269 19558 50303
rect 21373 50269 21407 50303
rect 22661 50269 22695 50303
rect 22753 50269 22787 50303
rect 22845 50269 22879 50303
rect 23029 50269 23063 50303
rect 23581 50269 23615 50303
rect 27813 50269 27847 50303
rect 29929 50269 29963 50303
rect 30205 50269 30239 50303
rect 32321 50269 32355 50303
rect 33241 50269 33275 50303
rect 35173 50269 35207 50303
rect 36093 50269 36127 50303
rect 36369 50269 36403 50303
rect 38301 50269 38335 50303
rect 38577 50269 38611 50303
rect 38761 50269 38795 50303
rect 39957 50269 39991 50303
rect 41245 50269 41279 50303
rect 45845 50269 45879 50303
rect 47041 50269 47075 50303
rect 47317 50269 47351 50303
rect 48145 50269 48179 50303
rect 48513 50269 48547 50303
rect 48881 50269 48915 50303
rect 50353 50269 50387 50303
rect 50537 50269 50571 50303
rect 51549 50269 51583 50303
rect 51816 50269 51850 50303
rect 23857 50201 23891 50235
rect 24593 50201 24627 50235
rect 26249 50201 26283 50235
rect 37565 50201 37599 50235
rect 38669 50201 38703 50235
rect 46213 50201 46247 50235
rect 12633 50133 12667 50167
rect 15393 50133 15427 50167
rect 16865 50133 16899 50167
rect 20637 50133 20671 50167
rect 22385 50133 22419 50167
rect 33425 50133 33459 50167
rect 35449 50133 35483 50167
rect 37657 50133 37691 50167
rect 40141 50133 40175 50167
rect 45937 50133 45971 50167
rect 46029 50133 46063 50167
rect 47501 50133 47535 50167
rect 48145 50133 48179 50167
rect 20269 49929 20303 49963
rect 24961 49929 24995 49963
rect 33517 49929 33551 49963
rect 36645 49929 36679 49963
rect 37473 49929 37507 49963
rect 43729 49929 43763 49963
rect 46489 49929 46523 49963
rect 49157 49929 49191 49963
rect 50537 49929 50571 49963
rect 51365 49929 51399 49963
rect 19901 49861 19935 49895
rect 20101 49861 20135 49895
rect 34621 49861 34655 49895
rect 35265 49861 35299 49895
rect 38301 49861 38335 49895
rect 41688 49861 41722 49895
rect 43361 49861 43395 49895
rect 43545 49861 43579 49895
rect 44833 49861 44867 49895
rect 48145 49861 48179 49895
rect 50077 49861 50111 49895
rect 12449 49793 12483 49827
rect 12716 49793 12750 49827
rect 14289 49793 14323 49827
rect 14545 49793 14579 49827
rect 16865 49793 16899 49827
rect 18638 49793 18672 49827
rect 24777 49793 24811 49827
rect 26249 49793 26283 49827
rect 28825 49793 28859 49827
rect 29377 49793 29411 49827
rect 30205 49793 30239 49827
rect 30472 49793 30506 49827
rect 32137 49793 32171 49827
rect 32404 49793 32438 49827
rect 34253 49793 34287 49827
rect 35449 49793 35483 49827
rect 35633 49793 35667 49827
rect 35725 49793 35759 49827
rect 36553 49793 36587 49827
rect 37381 49793 37415 49827
rect 38485 49793 38519 49827
rect 39497 49793 39531 49827
rect 39957 49793 39991 49827
rect 42441 49793 42475 49827
rect 44741 49793 44775 49827
rect 44925 49793 44959 49827
rect 45043 49793 45077 49827
rect 45937 49793 45971 49827
rect 48789 49793 48823 49827
rect 50353 49793 50387 49827
rect 51273 49793 51307 49827
rect 52101 49793 52135 49827
rect 17601 49725 17635 49759
rect 17785 49725 17819 49759
rect 18521 49725 18555 49759
rect 18797 49725 18831 49759
rect 19441 49725 19475 49759
rect 22477 49725 22511 49759
rect 22661 49725 22695 49759
rect 23857 49725 23891 49759
rect 29653 49725 29687 49759
rect 40325 49725 40359 49759
rect 44557 49725 44591 49759
rect 45201 49725 45235 49759
rect 46213 49725 46247 49759
rect 47777 49725 47811 49759
rect 48881 49725 48915 49759
rect 50261 49725 50295 49759
rect 13829 49657 13863 49691
rect 15669 49657 15703 49691
rect 18245 49657 18279 49691
rect 31585 49657 31619 49691
rect 39405 49657 39439 49691
rect 41889 49657 41923 49691
rect 48329 49657 48363 49691
rect 16865 49589 16899 49623
rect 20085 49589 20119 49623
rect 26065 49589 26099 49623
rect 28641 49589 28675 49623
rect 34621 49589 34655 49623
rect 34805 49589 34839 49623
rect 42625 49589 42659 49623
rect 43545 49589 43579 49623
rect 46305 49589 46339 49623
rect 48145 49589 48179 49623
rect 48973 49589 49007 49623
rect 50077 49589 50111 49623
rect 51917 49589 51951 49623
rect 14381 49385 14415 49419
rect 17693 49385 17727 49419
rect 18521 49385 18555 49419
rect 19349 49385 19383 49419
rect 23029 49385 23063 49419
rect 31125 49385 31159 49419
rect 36093 49385 36127 49419
rect 39129 49385 39163 49419
rect 46305 49385 46339 49419
rect 48789 49385 48823 49419
rect 51273 49385 51307 49419
rect 40141 49317 40175 49351
rect 13093 49249 13127 49283
rect 18153 49249 18187 49283
rect 20177 49249 20211 49283
rect 38393 49249 38427 49283
rect 40877 49249 40911 49283
rect 13277 49181 13311 49215
rect 14565 49181 14599 49215
rect 15025 49181 15059 49215
rect 15301 49181 15335 49215
rect 16313 49181 16347 49215
rect 18337 49181 18371 49215
rect 19257 49181 19291 49215
rect 19901 49181 19935 49215
rect 21649 49181 21683 49215
rect 24869 49181 24903 49215
rect 24961 49181 24995 49215
rect 25513 49181 25547 49215
rect 25780 49181 25814 49215
rect 27629 49181 27663 49215
rect 27896 49181 27930 49215
rect 30297 49181 30331 49215
rect 31309 49181 31343 49215
rect 32597 49181 32631 49215
rect 34713 49181 34747 49215
rect 37105 49181 37139 49215
rect 38301 49181 38335 49215
rect 38945 49181 38979 49215
rect 39865 49181 39899 49215
rect 40601 49181 40635 49215
rect 41429 49181 41463 49215
rect 41613 49181 41647 49215
rect 41981 49181 42015 49215
rect 43453 49181 43487 49215
rect 43729 49181 43763 49215
rect 43913 49181 43947 49215
rect 45201 49181 45235 49215
rect 45385 49181 45419 49215
rect 45661 49181 45695 49215
rect 46121 49181 46155 49215
rect 46489 49181 46523 49215
rect 48697 49181 48731 49215
rect 49341 49181 49375 49215
rect 49525 49181 49559 49215
rect 50997 49181 51031 49215
rect 51089 49181 51123 49215
rect 51733 49181 51767 49215
rect 52000 49181 52034 49215
rect 16580 49113 16614 49147
rect 21916 49113 21950 49147
rect 30665 49113 30699 49147
rect 32965 49113 32999 49147
rect 33609 49113 33643 49147
rect 34958 49113 34992 49147
rect 42901 49113 42935 49147
rect 45017 49113 45051 49147
rect 45293 49113 45327 49147
rect 45503 49113 45537 49147
rect 49433 49113 49467 49147
rect 13461 49045 13495 49079
rect 26893 49045 26927 49079
rect 29009 49045 29043 49079
rect 33701 49045 33735 49079
rect 37289 49045 37323 49079
rect 41613 49045 41647 49079
rect 46673 49045 46707 49079
rect 53113 49045 53147 49079
rect 13001 48841 13035 48875
rect 19625 48841 19659 48875
rect 21189 48841 21223 48875
rect 26341 48841 26375 48875
rect 27353 48841 27387 48875
rect 29469 48841 29503 48875
rect 34621 48841 34655 48875
rect 36553 48841 36587 48875
rect 41705 48841 41739 48875
rect 43913 48841 43947 48875
rect 45937 48841 45971 48875
rect 46029 48841 46063 48875
rect 46949 48841 46983 48875
rect 47803 48841 47837 48875
rect 51641 48841 51675 48875
rect 17325 48773 17359 48807
rect 29101 48773 29135 48807
rect 29301 48773 29335 48807
rect 30021 48773 30055 48807
rect 37534 48773 37568 48807
rect 45845 48773 45879 48807
rect 47593 48773 47627 48807
rect 50537 48773 50571 48807
rect 13185 48705 13219 48739
rect 14013 48705 14047 48739
rect 17141 48705 17175 48739
rect 19809 48705 19843 48739
rect 20269 48705 20303 48739
rect 21005 48705 21039 48739
rect 24777 48705 24811 48739
rect 24961 48705 24995 48739
rect 25605 48705 25639 48739
rect 26249 48705 26283 48739
rect 27169 48705 27203 48739
rect 28825 48705 28859 48739
rect 34805 48705 34839 48739
rect 36737 48705 36771 48739
rect 39865 48705 39899 48739
rect 39957 48705 39991 48739
rect 40693 48705 40727 48739
rect 41521 48705 41555 48739
rect 42993 48705 43027 48739
rect 43729 48705 43763 48739
rect 43913 48705 43947 48739
rect 46213 48705 46247 48739
rect 46765 48705 46799 48739
rect 47041 48705 47075 48739
rect 48881 48705 48915 48739
rect 49617 48705 49651 48739
rect 50353 48705 50387 48739
rect 51457 48705 51491 48739
rect 24593 48637 24627 48671
rect 26985 48637 27019 48671
rect 37289 48637 37323 48671
rect 40141 48637 40175 48671
rect 41337 48637 41371 48671
rect 42809 48637 42843 48671
rect 43085 48637 43119 48671
rect 43177 48637 43211 48671
rect 30205 48569 30239 48603
rect 40049 48569 40083 48603
rect 45661 48569 45695 48603
rect 14197 48501 14231 48535
rect 20453 48501 20487 48535
rect 25421 48501 25455 48535
rect 29285 48501 29319 48535
rect 38669 48501 38703 48535
rect 40785 48501 40819 48535
rect 46765 48501 46799 48535
rect 47777 48501 47811 48535
rect 47961 48501 47995 48535
rect 48973 48501 49007 48535
rect 49709 48501 49743 48535
rect 19809 48297 19843 48331
rect 19993 48297 20027 48331
rect 41613 48297 41647 48331
rect 43821 48297 43855 48331
rect 45385 48297 45419 48331
rect 45845 48297 45879 48331
rect 32229 48229 32263 48263
rect 32873 48229 32907 48263
rect 37381 48229 37415 48263
rect 41797 48229 41831 48263
rect 43085 48229 43119 48263
rect 47041 48229 47075 48263
rect 49249 48229 49283 48263
rect 20453 48161 20487 48195
rect 33701 48161 33735 48195
rect 33885 48161 33919 48195
rect 40325 48161 40359 48195
rect 43545 48161 43579 48195
rect 44373 48161 44407 48195
rect 45569 48161 45603 48195
rect 47225 48161 47259 48195
rect 50169 48161 50203 48195
rect 1961 48093 1995 48127
rect 12909 48093 12943 48127
rect 14473 48093 14507 48127
rect 15209 48093 15243 48127
rect 15669 48093 15703 48127
rect 16497 48093 16531 48127
rect 17233 48093 17267 48127
rect 20720 48093 20754 48127
rect 23213 48093 23247 48127
rect 23305 48093 23339 48127
rect 24409 48093 24443 48127
rect 24676 48093 24710 48127
rect 26341 48093 26375 48127
rect 27353 48093 27387 48127
rect 29745 48093 29779 48127
rect 30481 48093 30515 48127
rect 31309 48093 31343 48127
rect 33149 48093 33183 48127
rect 33609 48093 33643 48127
rect 37105 48093 37139 48127
rect 37197 48093 37231 48127
rect 40049 48093 40083 48127
rect 40233 48093 40267 48127
rect 44281 48093 44315 48127
rect 44465 48093 44499 48127
rect 45293 48093 45327 48127
rect 46949 48093 46983 48127
rect 48513 48093 48547 48127
rect 48789 48093 48823 48127
rect 49433 48093 49467 48127
rect 49525 48093 49559 48127
rect 50425 48093 50459 48127
rect 15761 48025 15795 48059
rect 19625 48025 19659 48059
rect 32045 48025 32079 48059
rect 32873 48025 32907 48059
rect 33885 48025 33919 48059
rect 41429 48025 41463 48059
rect 41629 48025 41663 48059
rect 43085 48025 43119 48059
rect 48329 48025 48363 48059
rect 49249 48025 49283 48059
rect 67741 48025 67775 48059
rect 12725 47957 12759 47991
rect 14473 47957 14507 47991
rect 15025 47957 15059 47991
rect 16497 47957 16531 47991
rect 17049 47957 17083 47991
rect 19835 47957 19869 47991
rect 21833 47957 21867 47991
rect 23489 47957 23523 47991
rect 25789 47957 25823 47991
rect 26433 47957 26467 47991
rect 27169 47957 27203 47991
rect 29837 47957 29871 47991
rect 30573 47957 30607 47991
rect 31125 47957 31159 47991
rect 33057 47957 33091 47991
rect 39865 47957 39899 47991
rect 43637 47957 43671 47991
rect 47225 47957 47259 47991
rect 48697 47957 48731 47991
rect 51549 47957 51583 47991
rect 67833 47957 67867 47991
rect 17417 47753 17451 47787
rect 24317 47753 24351 47787
rect 27537 47753 27571 47787
rect 34989 47753 35023 47787
rect 35817 47753 35851 47787
rect 12440 47685 12474 47719
rect 14464 47685 14498 47719
rect 28181 47685 28215 47719
rect 28549 47685 28583 47719
rect 28917 47685 28951 47719
rect 29285 47685 29319 47719
rect 30472 47685 30506 47719
rect 36093 47685 36127 47719
rect 40877 47685 40911 47719
rect 43269 47685 43303 47719
rect 48329 47685 48363 47719
rect 48697 47685 48731 47719
rect 1685 47617 1719 47651
rect 14197 47617 14231 47651
rect 17233 47617 17267 47651
rect 18061 47617 18095 47651
rect 22293 47617 22327 47651
rect 22560 47617 22594 47651
rect 24317 47617 24351 47651
rect 26249 47617 26283 47651
rect 27261 47617 27295 47651
rect 27353 47617 27387 47651
rect 28457 47617 28491 47651
rect 30205 47617 30239 47651
rect 32597 47617 32631 47651
rect 32864 47617 32898 47651
rect 34805 47617 34839 47651
rect 35081 47617 35115 47651
rect 35725 47617 35759 47651
rect 35909 47617 35943 47651
rect 37841 47617 37875 47651
rect 39037 47617 39071 47651
rect 39405 47617 39439 47651
rect 39773 47617 39807 47651
rect 40693 47617 40727 47651
rect 40969 47617 41003 47651
rect 41429 47617 41463 47651
rect 41613 47617 41647 47651
rect 43729 47617 43763 47651
rect 44925 47617 44959 47651
rect 45201 47617 45235 47651
rect 48513 47617 48547 47651
rect 50353 47617 50387 47651
rect 50445 47617 50479 47651
rect 50629 47617 50663 47651
rect 50721 47617 50755 47651
rect 51641 47617 51675 47651
rect 1869 47549 1903 47583
rect 2789 47549 2823 47583
rect 12173 47549 12207 47583
rect 17049 47549 17083 47583
rect 17877 47549 17911 47583
rect 18797 47549 18831 47583
rect 18914 47549 18948 47583
rect 19073 47549 19107 47583
rect 39865 47549 39899 47583
rect 43637 47549 43671 47583
rect 45109 47549 45143 47583
rect 50169 47549 50203 47583
rect 15577 47481 15611 47515
rect 18521 47481 18555 47515
rect 35541 47481 35575 47515
rect 40141 47481 40175 47515
rect 43913 47481 43947 47515
rect 45385 47481 45419 47515
rect 13553 47413 13587 47447
rect 19717 47413 19751 47447
rect 23673 47413 23707 47447
rect 26341 47413 26375 47447
rect 29469 47413 29503 47447
rect 31585 47413 31619 47447
rect 33977 47413 34011 47447
rect 34621 47413 34655 47447
rect 38025 47413 38059 47447
rect 40693 47413 40727 47447
rect 41429 47413 41463 47447
rect 43361 47413 43395 47447
rect 45201 47413 45235 47447
rect 51457 47413 51491 47447
rect 2421 47209 2455 47243
rect 12265 47209 12299 47243
rect 13369 47209 13403 47243
rect 15301 47209 15335 47243
rect 17693 47209 17727 47243
rect 23121 47209 23155 47243
rect 27813 47209 27847 47243
rect 30389 47209 30423 47243
rect 30573 47209 30607 47243
rect 33977 47209 34011 47243
rect 40049 47209 40083 47243
rect 40233 47209 40267 47243
rect 45385 47209 45419 47243
rect 45845 47209 45879 47243
rect 46305 47209 46339 47243
rect 46673 47209 46707 47243
rect 53021 47209 53055 47243
rect 29929 47141 29963 47175
rect 34161 47141 34195 47175
rect 34989 47141 35023 47175
rect 41245 47141 41279 47175
rect 13001 47073 13035 47107
rect 14933 47073 14967 47107
rect 16313 47073 16347 47107
rect 22109 47073 22143 47107
rect 26433 47073 26467 47107
rect 40785 47073 40819 47107
rect 45569 47073 45603 47107
rect 2329 47005 2363 47039
rect 12357 47005 12391 47039
rect 13185 47005 13219 47039
rect 15117 47005 15151 47039
rect 16580 47005 16614 47039
rect 20269 47005 20303 47039
rect 21005 47005 21039 47039
rect 21833 47005 21867 47039
rect 23305 47005 23339 47039
rect 26700 47005 26734 47039
rect 28733 47005 28767 47039
rect 31677 47005 31711 47039
rect 32505 47005 32539 47039
rect 35725 47005 35759 47039
rect 36093 47005 36127 47039
rect 36461 47005 36495 47039
rect 36737 47005 36771 47039
rect 37657 47005 37691 47039
rect 38025 47005 38059 47039
rect 38209 47005 38243 47039
rect 38945 47005 38979 47039
rect 40877 47005 40911 47039
rect 44189 47005 44223 47039
rect 45385 47005 45419 47039
rect 45661 47005 45695 47039
rect 46305 47005 46339 47039
rect 46397 47005 46431 47039
rect 50997 47005 51031 47039
rect 51181 47005 51215 47039
rect 51641 47005 51675 47039
rect 51897 47005 51931 47039
rect 67925 47005 67959 47039
rect 30205 46937 30239 46971
rect 30405 46937 30439 46971
rect 33793 46937 33827 46971
rect 34009 46937 34043 46971
rect 34805 46937 34839 46971
rect 36645 46937 36679 46971
rect 39865 46937 39899 46971
rect 40065 46937 40099 46971
rect 44005 46937 44039 46971
rect 20269 46869 20303 46903
rect 20821 46869 20855 46903
rect 28917 46869 28951 46903
rect 31861 46869 31895 46903
rect 32597 46869 32631 46903
rect 37473 46869 37507 46903
rect 36461 46665 36495 46699
rect 42625 46665 42659 46699
rect 43177 46665 43211 46699
rect 45845 46665 45879 46699
rect 48973 46665 49007 46699
rect 50813 46665 50847 46699
rect 51917 46665 51951 46699
rect 20168 46597 20202 46631
rect 34069 46597 34103 46631
rect 47838 46597 47872 46631
rect 49700 46597 49734 46631
rect 1869 46529 1903 46563
rect 17417 46529 17451 46563
rect 17509 46529 17543 46563
rect 19073 46529 19107 46563
rect 19901 46529 19935 46563
rect 21833 46529 21867 46563
rect 22753 46529 22787 46563
rect 24041 46529 24075 46563
rect 24961 46529 24995 46563
rect 28549 46529 28583 46563
rect 29285 46529 29319 46563
rect 30021 46529 30055 46563
rect 30941 46529 30975 46563
rect 36369 46529 36403 46563
rect 37749 46529 37783 46563
rect 38577 46529 38611 46563
rect 39405 46529 39439 46563
rect 39497 46529 39531 46563
rect 41705 46529 41739 46563
rect 41889 46529 41923 46563
rect 42533 46529 42567 46563
rect 43361 46529 43395 46563
rect 43637 46529 43671 46563
rect 44465 46529 44499 46563
rect 45477 46529 45511 46563
rect 45661 46529 45695 46563
rect 46949 46529 46983 46563
rect 51549 46529 51583 46563
rect 51733 46529 51767 46563
rect 65809 46529 65843 46563
rect 24225 46461 24259 46495
rect 25078 46461 25112 46495
rect 25237 46461 25271 46495
rect 32781 46461 32815 46495
rect 33057 46461 33091 46495
rect 35817 46461 35851 46495
rect 39681 46461 39715 46495
rect 44189 46461 44223 46495
rect 47041 46461 47075 46495
rect 47593 46461 47627 46495
rect 49433 46461 49467 46495
rect 65993 46461 66027 46495
rect 67557 46461 67591 46495
rect 2053 46393 2087 46427
rect 24685 46393 24719 46427
rect 38025 46393 38059 46427
rect 43453 46393 43487 46427
rect 43545 46393 43579 46427
rect 17693 46325 17727 46359
rect 19257 46325 19291 46359
rect 21281 46325 21315 46359
rect 21833 46325 21867 46359
rect 22569 46325 22603 46359
rect 25881 46325 25915 46359
rect 28641 46325 28675 46359
rect 29469 46325 29503 46359
rect 30021 46325 30055 46359
rect 30757 46325 30791 46359
rect 38761 46325 38795 46359
rect 39589 46325 39623 46359
rect 41797 46325 41831 46359
rect 45477 46325 45511 46359
rect 17877 46121 17911 46155
rect 19901 46121 19935 46155
rect 20729 46121 20763 46155
rect 35081 46121 35115 46155
rect 36829 46121 36863 46155
rect 41429 46121 41463 46155
rect 43453 46121 43487 46155
rect 45201 46121 45235 46155
rect 45845 46121 45879 46155
rect 48237 46121 48271 46155
rect 67373 46121 67407 46155
rect 20085 46053 20119 46087
rect 45109 46053 45143 46087
rect 21649 45985 21683 46019
rect 24777 45985 24811 46019
rect 29929 45985 29963 46019
rect 32045 45985 32079 46019
rect 50629 45985 50663 46019
rect 13185 45917 13219 45951
rect 14473 45917 14507 45951
rect 15393 45917 15427 45951
rect 16497 45917 16531 45951
rect 18521 45917 18555 45951
rect 21916 45917 21950 45951
rect 23857 45917 23891 45951
rect 24501 45917 24535 45951
rect 24593 45917 24627 45951
rect 25789 45917 25823 45951
rect 28549 45917 28583 45951
rect 30196 45917 30230 45951
rect 34069 45917 34103 45951
rect 34713 45917 34747 45951
rect 35817 45917 35851 45951
rect 40049 45917 40083 45951
rect 40305 45917 40339 45951
rect 42073 45917 42107 45951
rect 42329 45917 42363 45951
rect 45017 45917 45051 45951
rect 45293 45917 45327 45951
rect 45753 45917 45787 45951
rect 48053 45917 48087 45951
rect 50813 45917 50847 45951
rect 50997 45917 51031 45951
rect 51641 45917 51675 45951
rect 67281 45917 67315 45951
rect 16764 45849 16798 45883
rect 19717 45849 19751 45883
rect 19933 45849 19967 45883
rect 20545 45849 20579 45883
rect 26034 45849 26068 45883
rect 32312 45849 32346 45883
rect 35081 45849 35115 45883
rect 36737 45849 36771 45883
rect 13001 45781 13035 45815
rect 14657 45781 14691 45815
rect 15209 45781 15243 45815
rect 18337 45781 18371 45815
rect 20745 45781 20779 45815
rect 20913 45781 20947 45815
rect 23029 45781 23063 45815
rect 23673 45781 23707 45815
rect 27169 45781 27203 45815
rect 28365 45781 28399 45815
rect 31309 45781 31343 45815
rect 33425 45781 33459 45815
rect 33885 45781 33919 45815
rect 35265 45781 35299 45815
rect 36093 45781 36127 45815
rect 51457 45781 51491 45815
rect 16865 45577 16899 45611
rect 22293 45577 22327 45611
rect 24685 45577 24719 45611
rect 29837 45577 29871 45611
rect 30757 45577 30791 45611
rect 42625 45577 42659 45611
rect 45385 45577 45419 45611
rect 12808 45509 12842 45543
rect 14832 45509 14866 45543
rect 19349 45509 19383 45543
rect 21925 45509 21959 45543
rect 22125 45509 22159 45543
rect 23572 45509 23606 45543
rect 25605 45509 25639 45543
rect 25805 45509 25839 45543
rect 27896 45509 27930 45543
rect 29469 45509 29503 45543
rect 29685 45509 29719 45543
rect 30389 45509 30423 45543
rect 30605 45509 30639 45543
rect 32689 45509 32723 45543
rect 32905 45509 32939 45543
rect 39396 45509 39430 45543
rect 50436 45509 50470 45543
rect 1869 45441 1903 45475
rect 14565 45441 14599 45475
rect 16865 45441 16899 45475
rect 17509 45441 17543 45475
rect 17693 45441 17727 45475
rect 18429 45441 18463 45475
rect 20076 45441 20110 45475
rect 26985 45441 27019 45475
rect 34161 45441 34195 45475
rect 35633 45441 35667 45475
rect 36461 45441 36495 45475
rect 37289 45441 37323 45475
rect 37556 45441 37590 45475
rect 41153 45441 41187 45475
rect 42441 45441 42475 45475
rect 44925 45441 44959 45475
rect 45201 45441 45235 45475
rect 47777 45441 47811 45475
rect 48513 45441 48547 45475
rect 12541 45373 12575 45407
rect 18546 45373 18580 45407
rect 18705 45373 18739 45407
rect 19809 45373 19843 45407
rect 23305 45373 23339 45407
rect 27077 45373 27111 45407
rect 27629 45373 27663 45407
rect 34437 45373 34471 45407
rect 36645 45373 36679 45407
rect 36737 45373 36771 45407
rect 39129 45373 39163 45407
rect 45109 45373 45143 45407
rect 50169 45373 50203 45407
rect 18153 45305 18187 45339
rect 33057 45305 33091 45339
rect 40509 45305 40543 45339
rect 1961 45237 1995 45271
rect 13921 45237 13955 45271
rect 15945 45237 15979 45271
rect 21189 45237 21223 45271
rect 22109 45237 22143 45271
rect 25789 45237 25823 45271
rect 25973 45237 26007 45271
rect 29009 45237 29043 45271
rect 29653 45237 29687 45271
rect 30573 45237 30607 45271
rect 32873 45237 32907 45271
rect 35449 45237 35483 45271
rect 36277 45237 36311 45271
rect 38669 45237 38703 45271
rect 40969 45237 41003 45271
rect 45201 45237 45235 45271
rect 47593 45237 47627 45271
rect 48329 45237 48363 45271
rect 51549 45237 51583 45271
rect 67649 45237 67683 45271
rect 12633 45033 12667 45067
rect 13553 45033 13587 45067
rect 15485 45033 15519 45067
rect 19441 45033 19475 45067
rect 19993 45033 20027 45067
rect 21465 45033 21499 45067
rect 25789 45033 25823 45067
rect 27629 45033 27663 45067
rect 28917 45033 28951 45067
rect 37473 45033 37507 45067
rect 40141 45033 40175 45067
rect 45477 45033 45511 45067
rect 50169 45033 50203 45067
rect 30481 44965 30515 44999
rect 45661 44965 45695 44999
rect 13185 44897 13219 44931
rect 15117 44897 15151 44931
rect 34897 44897 34931 44931
rect 38117 44897 38151 44931
rect 45385 44897 45419 44931
rect 47593 44897 47627 44931
rect 66269 44897 66303 44931
rect 68109 44897 68143 44931
rect 12633 44829 12667 44863
rect 13369 44829 13403 44863
rect 15301 44829 15335 44863
rect 19441 44829 19475 44863
rect 20177 44829 20211 44863
rect 21649 44829 21683 44863
rect 21925 44829 21959 44863
rect 23029 44829 23063 44863
rect 25973 44829 26007 44863
rect 27537 44829 27571 44863
rect 28733 44829 28767 44863
rect 31125 44829 31159 44863
rect 32505 44829 32539 44863
rect 35164 44829 35198 44863
rect 37657 44829 37691 44863
rect 38301 44829 38335 44863
rect 40141 44829 40175 44863
rect 41705 44829 41739 44863
rect 41961 44829 41995 44863
rect 44005 44829 44039 44863
rect 45477 44829 45511 44863
rect 46305 44829 46339 44863
rect 47860 44829 47894 44863
rect 50353 44829 50387 44863
rect 23121 44761 23155 44795
rect 30297 44761 30331 44795
rect 38485 44761 38519 44795
rect 45017 44761 45051 44795
rect 66453 44761 66487 44795
rect 21833 44693 21867 44727
rect 31125 44693 31159 44727
rect 32597 44693 32631 44727
rect 36277 44693 36311 44727
rect 43085 44693 43119 44727
rect 43821 44693 43855 44727
rect 46535 44693 46569 44727
rect 48973 44693 49007 44727
rect 14657 44489 14691 44523
rect 23397 44489 23431 44523
rect 30957 44489 30991 44523
rect 31125 44489 31159 44523
rect 34805 44489 34839 44523
rect 41797 44489 41831 44523
rect 44557 44489 44591 44523
rect 45845 44489 45879 44523
rect 47961 44489 47995 44523
rect 49433 44489 49467 44523
rect 67557 44489 67591 44523
rect 22753 44421 22787 44455
rect 30757 44421 30791 44455
rect 35624 44421 35658 44455
rect 12633 44353 12667 44387
rect 14473 44353 14507 44387
rect 15393 44353 15427 44387
rect 16865 44353 16899 44387
rect 18153 44353 18187 44387
rect 22569 44353 22603 44387
rect 22845 44353 22879 44387
rect 23305 44353 23339 44387
rect 25237 44353 25271 44387
rect 27169 44353 27203 44387
rect 30113 44353 30147 44387
rect 32321 44353 32355 44387
rect 33977 44353 34011 44387
rect 34713 44353 34747 44387
rect 35357 44353 35391 44387
rect 41613 44353 41647 44387
rect 42441 44353 42475 44387
rect 43444 44353 43478 44387
rect 45477 44353 45511 44387
rect 46305 44353 46339 44387
rect 47685 44353 47719 44387
rect 47777 44353 47811 44387
rect 48513 44353 48547 44387
rect 49249 44353 49283 44387
rect 67465 44353 67499 44387
rect 17969 44285 18003 44319
rect 18889 44285 18923 44319
rect 19006 44285 19040 44319
rect 19165 44285 19199 44319
rect 43177 44285 43211 44319
rect 45569 44285 45603 44319
rect 18613 44217 18647 44251
rect 42625 44217 42659 44251
rect 46397 44217 46431 44251
rect 12633 44149 12667 44183
rect 15209 44149 15243 44183
rect 16681 44149 16715 44183
rect 19809 44149 19843 44183
rect 22385 44149 22419 44183
rect 25053 44149 25087 44183
rect 26985 44149 27019 44183
rect 30205 44149 30239 44183
rect 30941 44149 30975 44183
rect 32137 44149 32171 44183
rect 33793 44149 33827 44183
rect 36737 44149 36771 44183
rect 45477 44149 45511 44183
rect 48605 44149 48639 44183
rect 1961 43945 1995 43979
rect 29745 43945 29779 43979
rect 36461 43945 36495 43979
rect 40233 43945 40267 43979
rect 42533 43945 42567 43979
rect 44373 43945 44407 43979
rect 16037 43877 16071 43911
rect 20361 43877 20395 43911
rect 25789 43877 25823 43911
rect 27813 43877 27847 43911
rect 29929 43877 29963 43911
rect 27353 43809 27387 43843
rect 28206 43809 28240 43843
rect 30941 43809 30975 43843
rect 36553 43809 36587 43843
rect 44005 43809 44039 43843
rect 45661 43809 45695 43843
rect 66269 43809 66303 43843
rect 13277 43741 13311 43775
rect 13369 43741 13403 43775
rect 14657 43741 14691 43775
rect 14924 43741 14958 43775
rect 16773 43741 16807 43775
rect 17029 43741 17063 43775
rect 20177 43741 20211 43775
rect 21097 43741 21131 43775
rect 21373 43741 21407 43775
rect 22017 43741 22051 43775
rect 22293 43741 22327 43775
rect 22753 43741 22787 43775
rect 23029 43741 23063 43775
rect 24409 43741 24443 43775
rect 24676 43741 24710 43775
rect 26249 43741 26283 43775
rect 27169 43741 27203 43775
rect 28089 43741 28123 43775
rect 28365 43741 28399 43775
rect 29009 43741 29043 43775
rect 31208 43741 31242 43775
rect 32781 43741 32815 43775
rect 33048 43741 33082 43775
rect 36277 43741 36311 43775
rect 37933 43741 37967 43775
rect 38117 43741 38151 43775
rect 38209 43741 38243 43775
rect 40049 43741 40083 43775
rect 40877 43741 40911 43775
rect 42441 43741 42475 43775
rect 44189 43741 44223 43775
rect 48053 43741 48087 43775
rect 1869 43673 1903 43707
rect 22201 43673 22235 43707
rect 29561 43673 29595 43707
rect 29777 43673 29811 43707
rect 36093 43673 36127 43707
rect 38669 43673 38703 43707
rect 38853 43673 38887 43707
rect 41061 43673 41095 43707
rect 45928 43673 45962 43707
rect 48320 43673 48354 43707
rect 66453 43673 66487 43707
rect 68109 43673 68143 43707
rect 13553 43605 13587 43639
rect 18153 43605 18187 43639
rect 20913 43605 20947 43639
rect 21281 43605 21315 43639
rect 21833 43605 21867 43639
rect 26433 43605 26467 43639
rect 32321 43605 32355 43639
rect 34161 43605 34195 43639
rect 39037 43605 39071 43639
rect 47041 43605 47075 43639
rect 49433 43605 49467 43639
rect 14749 43401 14783 43435
rect 15669 43401 15703 43435
rect 17049 43401 17083 43435
rect 24133 43401 24167 43435
rect 25697 43401 25731 43435
rect 28365 43401 28399 43435
rect 33241 43401 33275 43435
rect 34161 43401 34195 43435
rect 40233 43401 40267 43435
rect 46397 43401 46431 43435
rect 48605 43401 48639 43435
rect 67557 43401 67591 43435
rect 27252 43333 27286 43367
rect 33793 43333 33827 43367
rect 33993 43333 34027 43367
rect 34713 43333 34747 43367
rect 38393 43333 38427 43367
rect 40785 43333 40819 43367
rect 12725 43265 12759 43299
rect 12992 43265 13026 43299
rect 14565 43265 14599 43299
rect 15393 43265 15427 43299
rect 15485 43265 15519 43299
rect 16773 43265 16807 43299
rect 16865 43265 16899 43299
rect 20294 43265 20328 43299
rect 22569 43265 22603 43299
rect 24041 43265 24075 43299
rect 25421 43265 25455 43299
rect 25513 43265 25547 43299
rect 26985 43265 27019 43299
rect 29377 43265 29411 43299
rect 33241 43265 33275 43299
rect 38025 43265 38059 43299
rect 39120 43265 39154 43299
rect 41797 43265 41831 43299
rect 44005 43265 44039 43299
rect 45661 43265 45695 43299
rect 45753 43265 45787 43299
rect 45937 43265 45971 43299
rect 46581 43265 46615 43299
rect 47685 43265 47719 43299
rect 47777 43265 47811 43299
rect 48421 43265 48455 43299
rect 67465 43265 67499 43299
rect 19257 43197 19291 43231
rect 19441 43197 19475 43231
rect 20177 43197 20211 43231
rect 20453 43197 20487 43231
rect 22845 43197 22879 43231
rect 29193 43197 29227 43231
rect 30113 43197 30147 43231
rect 30230 43197 30264 43231
rect 30389 43197 30423 43231
rect 38853 43197 38887 43231
rect 14105 43129 14139 43163
rect 19901 43129 19935 43163
rect 29837 43129 29871 43163
rect 40969 43129 41003 43163
rect 21097 43061 21131 43095
rect 31033 43061 31067 43095
rect 33977 43061 34011 43095
rect 34805 43061 34839 43095
rect 41797 43061 41831 43095
rect 43821 43061 43855 43095
rect 47961 43061 47995 43095
rect 13185 42857 13219 42891
rect 32597 42857 32631 42891
rect 33977 42857 34011 42891
rect 38945 42857 38979 42891
rect 32781 42789 32815 42823
rect 17601 42721 17635 42755
rect 36829 42721 36863 42755
rect 39865 42721 39899 42755
rect 44373 42721 44407 42755
rect 67925 42721 67959 42755
rect 13369 42653 13403 42687
rect 14749 42653 14783 42687
rect 15669 42653 15703 42687
rect 16957 42653 16991 42687
rect 17785 42653 17819 42687
rect 21373 42653 21407 42687
rect 21649 42653 21683 42687
rect 23673 42653 23707 42687
rect 23765 42653 23799 42687
rect 24409 42653 24443 42687
rect 29561 42653 29595 42687
rect 29837 42653 29871 42687
rect 30849 42653 30883 42687
rect 31953 42653 31987 42687
rect 34713 42653 34747 42687
rect 37105 42653 37139 42687
rect 38117 42653 38151 42687
rect 38301 42653 38335 42687
rect 38945 42653 38979 42687
rect 40049 42653 40083 42687
rect 41153 42653 41187 42687
rect 43177 42653 43211 42687
rect 45201 42653 45235 42687
rect 48145 42653 48179 42687
rect 67281 42653 67315 42687
rect 1869 42585 1903 42619
rect 21189 42585 21223 42619
rect 24654 42585 24688 42619
rect 32413 42585 32447 42619
rect 33793 42585 33827 42619
rect 34980 42585 35014 42619
rect 41420 42585 41454 42619
rect 44097 42585 44131 42619
rect 1961 42517 1995 42551
rect 14933 42517 14967 42551
rect 15485 42517 15519 42551
rect 17049 42517 17083 42551
rect 17969 42517 18003 42551
rect 21557 42517 21591 42551
rect 25789 42517 25823 42551
rect 31033 42517 31067 42551
rect 31769 42517 31803 42551
rect 32613 42517 32647 42551
rect 33993 42517 34027 42551
rect 34161 42517 34195 42551
rect 36093 42517 36127 42551
rect 38209 42517 38243 42551
rect 40233 42517 40267 42551
rect 42533 42517 42567 42551
rect 42993 42517 43027 42551
rect 45017 42517 45051 42551
rect 47961 42517 47995 42551
rect 18337 42313 18371 42347
rect 25605 42313 25639 42347
rect 28365 42313 28399 42347
rect 34161 42313 34195 42347
rect 35449 42313 35483 42347
rect 15016 42245 15050 42279
rect 22293 42245 22327 42279
rect 32382 42245 32416 42279
rect 34805 42245 34839 42279
rect 41613 42245 41647 42279
rect 43361 42245 43395 42279
rect 44088 42245 44122 42279
rect 14749 42177 14783 42211
rect 16957 42177 16991 42211
rect 17224 42177 17258 42211
rect 18797 42177 18831 42211
rect 19625 42177 19659 42211
rect 19717 42177 19751 42211
rect 22661 42177 22695 42211
rect 23213 42177 23247 42211
rect 23397 42177 23431 42211
rect 23857 42177 23891 42211
rect 24961 42177 24995 42211
rect 25053 42177 25087 42211
rect 25881 42177 25915 42211
rect 26157 42177 26191 42211
rect 26985 42177 27019 42211
rect 27445 42177 27479 42211
rect 27813 42177 27847 42211
rect 28365 42177 28399 42211
rect 29101 42177 29135 42211
rect 31309 42177 31343 42211
rect 33977 42177 34011 42211
rect 35633 42177 35667 42211
rect 36369 42177 36403 42211
rect 36553 42177 36587 42211
rect 37289 42177 37323 42211
rect 37473 42177 37507 42211
rect 38577 42177 38611 42211
rect 39773 42177 39807 42211
rect 41337 42177 41371 42211
rect 41429 42177 41463 42211
rect 43177 42177 43211 42211
rect 43821 42177 43855 42211
rect 65809 42177 65843 42211
rect 25973 42109 26007 42143
rect 31585 42109 31619 42143
rect 32126 42109 32160 42143
rect 38669 42109 38703 42143
rect 38761 42109 38795 42143
rect 38853 42109 38887 42143
rect 42993 42109 43027 42143
rect 48605 42109 48639 42143
rect 48789 42109 48823 42143
rect 50445 42109 50479 42143
rect 65993 42109 66027 42143
rect 67557 42109 67591 42143
rect 26341 42041 26375 42075
rect 36737 42041 36771 42075
rect 39589 42041 39623 42075
rect 16129 41973 16163 42007
rect 18981 41973 19015 42007
rect 19901 41973 19935 42007
rect 24041 41973 24075 42007
rect 25237 41973 25271 42007
rect 25881 41973 25915 42007
rect 28917 41973 28951 42007
rect 33517 41973 33551 42007
rect 34897 41973 34931 42007
rect 37657 41973 37691 42007
rect 38393 41973 38427 42007
rect 45201 41973 45235 42007
rect 15761 41769 15795 41803
rect 17049 41769 17083 41803
rect 17601 41769 17635 41803
rect 20637 41769 20671 41803
rect 23581 41769 23615 41803
rect 24409 41769 24443 41803
rect 25789 41769 25823 41803
rect 26433 41769 26467 41803
rect 26617 41769 26651 41803
rect 67649 41769 67683 41803
rect 17785 41701 17819 41735
rect 29009 41701 29043 41735
rect 49433 41701 49467 41735
rect 15393 41633 15427 41667
rect 17417 41633 17451 41667
rect 19257 41633 19291 41667
rect 26249 41633 26283 41667
rect 32321 41633 32355 41667
rect 41429 41633 41463 41667
rect 42246 41633 42280 41667
rect 42441 41633 42475 41667
rect 43361 41633 43395 41667
rect 15577 41565 15611 41599
rect 17601 41565 17635 41599
rect 21097 41565 21131 41599
rect 23397 41565 23431 41599
rect 24593 41565 24627 41599
rect 26157 41565 26191 41599
rect 26433 41565 26467 41599
rect 27629 41565 27663 41599
rect 29929 41565 29963 41599
rect 33241 41565 33275 41599
rect 35449 41565 35483 41599
rect 37197 41565 37231 41599
rect 37565 41565 37599 41599
rect 38623 41565 38657 41599
rect 38761 41565 38795 41599
rect 38858 41565 38892 41599
rect 39037 41565 39071 41599
rect 41245 41565 41279 41599
rect 42165 41565 42199 41599
rect 42349 41565 42383 41599
rect 43177 41565 43211 41599
rect 45477 41565 45511 41599
rect 45569 41565 45603 41599
rect 45661 41565 45695 41599
rect 45845 41565 45879 41599
rect 46305 41565 46339 41599
rect 48697 41565 48731 41599
rect 49341 41565 49375 41599
rect 67557 41565 67591 41599
rect 17325 41497 17359 41531
rect 19524 41497 19558 41531
rect 21364 41497 21398 41531
rect 27896 41497 27930 41531
rect 30196 41497 30230 41531
rect 32137 41497 32171 41531
rect 36553 41497 36587 41531
rect 37381 41497 37415 41531
rect 41061 41497 41095 41531
rect 42993 41497 43027 41531
rect 46550 41497 46584 41531
rect 22477 41429 22511 41463
rect 26985 41429 27019 41463
rect 31309 41429 31343 41463
rect 33333 41429 33367 41463
rect 35265 41429 35299 41463
rect 36645 41429 36679 41463
rect 38393 41429 38427 41463
rect 41981 41429 42015 41463
rect 45201 41429 45235 41463
rect 47685 41429 47719 41463
rect 48789 41429 48823 41463
rect 17417 41225 17451 41259
rect 19441 41225 19475 41259
rect 21833 41225 21867 41259
rect 23673 41225 23707 41259
rect 28733 41225 28767 41259
rect 29285 41225 29319 41259
rect 30665 41225 30699 41259
rect 42441 41225 42475 41259
rect 23397 41157 23431 41191
rect 27721 41157 27755 41191
rect 35164 41157 35198 41191
rect 39190 41157 39224 41191
rect 48881 41157 48915 41191
rect 17601 41089 17635 41123
rect 19625 41089 19659 41123
rect 22109 41089 22143 41123
rect 22201 41089 22235 41123
rect 22293 41089 22327 41123
rect 22477 41089 22511 41123
rect 24961 41089 24995 41123
rect 25421 41089 25455 41123
rect 27537 41089 27571 41123
rect 28457 41089 28491 41123
rect 28549 41089 28583 41123
rect 29193 41089 29227 41123
rect 30021 41089 30055 41123
rect 30205 41089 30239 41123
rect 30849 41089 30883 41123
rect 32505 41089 32539 41123
rect 32689 41089 32723 41123
rect 34897 41089 34931 41123
rect 37289 41089 37323 41123
rect 37473 41089 37507 41123
rect 38117 41089 38151 41123
rect 38945 41089 38979 41123
rect 42717 41089 42751 41123
rect 43453 41089 43487 41123
rect 44373 41089 44407 41123
rect 45983 41089 46017 41123
rect 46121 41089 46155 41123
rect 46213 41089 46247 41123
rect 46397 41089 46431 41123
rect 67465 41089 67499 41123
rect 29837 41021 29871 41055
rect 33425 41021 33459 41055
rect 33542 41021 33576 41055
rect 33701 41021 33735 41055
rect 41061 41021 41095 41055
rect 41337 41021 41371 41055
rect 42625 41021 42659 41055
rect 42809 41021 42843 41055
rect 42901 41021 42935 41055
rect 48697 41021 48731 41055
rect 50537 41021 50571 41055
rect 25513 40953 25547 40987
rect 33149 40953 33183 40987
rect 38301 40953 38335 40987
rect 24777 40885 24811 40919
rect 34345 40885 34379 40919
rect 36277 40885 36311 40919
rect 37657 40885 37691 40919
rect 40325 40885 40359 40919
rect 43637 40885 43671 40919
rect 44189 40885 44223 40919
rect 45753 40885 45787 40919
rect 67005 40885 67039 40919
rect 67557 40885 67591 40919
rect 35357 40681 35391 40715
rect 35541 40681 35575 40715
rect 36277 40681 36311 40715
rect 42901 40681 42935 40715
rect 43913 40681 43947 40715
rect 48053 40681 48087 40715
rect 27629 40613 27663 40647
rect 41061 40613 41095 40647
rect 19257 40545 19291 40579
rect 19717 40545 19751 40579
rect 24409 40545 24443 40579
rect 28089 40545 28123 40579
rect 38485 40545 38519 40579
rect 38577 40545 38611 40579
rect 38669 40545 38703 40579
rect 46673 40545 46707 40579
rect 66269 40545 66303 40579
rect 66453 40545 66487 40579
rect 68109 40545 68143 40579
rect 18521 40477 18555 40511
rect 21787 40477 21821 40511
rect 21925 40477 21959 40511
rect 22017 40477 22051 40511
rect 22201 40477 22235 40511
rect 23213 40477 23247 40511
rect 24676 40477 24710 40511
rect 26249 40477 26283 40511
rect 28273 40477 28307 40511
rect 29561 40477 29595 40511
rect 36461 40477 36495 40511
rect 38761 40477 38795 40511
rect 41245 40477 41279 40511
rect 43637 40477 43671 40511
rect 43729 40477 43763 40511
rect 45477 40477 45511 40511
rect 46929 40477 46963 40511
rect 48789 40477 48823 40511
rect 18613 40409 18647 40443
rect 19441 40409 19475 40443
rect 26516 40409 26550 40443
rect 35173 40409 35207 40443
rect 37013 40409 37047 40443
rect 42533 40409 42567 40443
rect 42717 40409 42751 40443
rect 21557 40341 21591 40375
rect 23397 40341 23431 40375
rect 25789 40341 25823 40375
rect 28457 40341 28491 40375
rect 29745 40341 29779 40375
rect 35373 40341 35407 40375
rect 37289 40341 37323 40375
rect 38301 40341 38335 40375
rect 45661 40341 45695 40375
rect 48881 40341 48915 40375
rect 25421 40137 25455 40171
rect 26341 40137 26375 40171
rect 26985 40137 27019 40171
rect 45201 40137 45235 40171
rect 32505 40069 32539 40103
rect 37289 40069 37323 40103
rect 38209 40069 38243 40103
rect 39037 40069 39071 40103
rect 42533 40069 42567 40103
rect 42717 40069 42751 40103
rect 48973 40069 49007 40103
rect 50629 40069 50663 40103
rect 67281 40069 67315 40103
rect 19901 40001 19935 40035
rect 20168 40001 20202 40035
rect 22661 40001 22695 40035
rect 22753 40001 22787 40035
rect 25145 40001 25179 40035
rect 25237 40001 25271 40035
rect 26341 40001 26375 40035
rect 27169 40001 27203 40035
rect 28273 40001 28307 40035
rect 29285 40001 29319 40035
rect 29552 40001 29586 40035
rect 31585 40001 31619 40035
rect 32321 40001 32355 40035
rect 33241 40001 33275 40035
rect 33425 40001 33459 40035
rect 35081 40001 35115 40035
rect 37473 40001 37507 40035
rect 40224 40001 40258 40035
rect 43821 40001 43855 40035
rect 44088 40001 44122 40035
rect 46351 40001 46385 40035
rect 46489 40001 46523 40035
rect 46581 40004 46615 40038
rect 46765 40001 46799 40035
rect 48789 40001 48823 40035
rect 27997 39933 28031 39967
rect 32137 39933 32171 39967
rect 34161 39933 34195 39967
rect 34278 39933 34312 39967
rect 34437 39933 34471 39967
rect 39957 39933 39991 39967
rect 33885 39865 33919 39899
rect 38393 39865 38427 39899
rect 1685 39797 1719 39831
rect 21281 39797 21315 39831
rect 30665 39797 30699 39831
rect 31401 39797 31435 39831
rect 37657 39797 37691 39831
rect 39129 39797 39163 39831
rect 41337 39797 41371 39831
rect 42901 39797 42935 39831
rect 46121 39797 46155 39831
rect 67373 39797 67407 39831
rect 25789 39593 25823 39627
rect 26525 39593 26559 39627
rect 30481 39593 30515 39627
rect 32689 39593 32723 39627
rect 35357 39593 35391 39627
rect 40233 39593 40267 39627
rect 42441 39593 42475 39627
rect 48145 39593 48179 39627
rect 1409 39457 1443 39491
rect 2789 39457 2823 39491
rect 19349 39457 19383 39491
rect 22477 39457 22511 39491
rect 29653 39457 29687 39491
rect 42717 39457 42751 39491
rect 42901 39457 42935 39491
rect 46765 39457 46799 39491
rect 26341 39389 26375 39423
rect 27261 39389 27295 39423
rect 28181 39389 28215 39423
rect 28273 39389 28307 39423
rect 29837 39389 29871 39423
rect 30021 39389 30055 39423
rect 30665 39389 30699 39423
rect 31309 39389 31343 39423
rect 31565 39389 31599 39423
rect 37473 39389 37507 39423
rect 38577 39389 38611 39423
rect 38666 39389 38700 39423
rect 38761 39389 38795 39423
rect 38945 39389 38979 39423
rect 40417 39389 40451 39423
rect 41061 39389 41095 39423
rect 41153 39389 41187 39423
rect 42625 39389 42659 39423
rect 42809 39389 42843 39423
rect 43637 39389 43671 39423
rect 45293 39389 45327 39423
rect 45382 39389 45416 39423
rect 45477 39383 45511 39417
rect 45661 39389 45695 39423
rect 46121 39389 46155 39423
rect 47021 39389 47055 39423
rect 48789 39389 48823 39423
rect 1593 39321 1627 39355
rect 19533 39321 19567 39355
rect 21189 39321 21223 39355
rect 22722 39321 22756 39355
rect 25513 39321 25547 39355
rect 35173 39321 35207 39355
rect 37289 39321 37323 39355
rect 37657 39321 37691 39355
rect 23857 39253 23891 39287
rect 27261 39253 27295 39287
rect 28457 39253 28491 39287
rect 35373 39253 35407 39287
rect 35541 39253 35575 39287
rect 38301 39253 38335 39287
rect 41337 39253 41371 39287
rect 43453 39253 43487 39287
rect 45017 39253 45051 39287
rect 46213 39253 46247 39287
rect 48881 39253 48915 39287
rect 1869 39049 1903 39083
rect 19717 39049 19751 39083
rect 22569 39049 22603 39083
rect 28457 39049 28491 39083
rect 31033 39049 31067 39083
rect 35265 39049 35299 39083
rect 39313 39049 39347 39083
rect 40509 39049 40543 39083
rect 42441 39049 42475 39083
rect 43821 39049 43855 39083
rect 46029 39049 46063 39083
rect 26433 38981 26467 39015
rect 41613 38981 41647 39015
rect 48973 38981 49007 39015
rect 1777 38913 1811 38947
rect 19625 38913 19659 38947
rect 20913 38913 20947 38947
rect 21005 38913 21039 38947
rect 21097 38913 21131 38947
rect 21281 38913 21315 38947
rect 22845 38913 22879 38947
rect 22937 38913 22971 38947
rect 23029 38913 23063 38947
rect 23213 38913 23247 38947
rect 23857 38913 23891 38947
rect 26249 38913 26283 38947
rect 27077 38913 27111 38947
rect 27344 38913 27378 38947
rect 30941 38913 30975 38947
rect 32321 38913 32355 38947
rect 33425 38913 33459 38947
rect 35817 38913 35851 38947
rect 36737 38913 36771 38947
rect 37933 38913 37967 38947
rect 38200 38913 38234 38947
rect 40693 38913 40727 38947
rect 41429 38913 41463 38947
rect 42717 38913 42751 38947
rect 42901 38913 42935 38947
rect 43453 38913 43487 38947
rect 43637 38913 43671 38947
rect 44649 38913 44683 38947
rect 44916 38913 44950 38947
rect 48789 38913 48823 38947
rect 24041 38845 24075 38879
rect 25605 38845 25639 38879
rect 32137 38845 32171 38879
rect 33609 38845 33643 38879
rect 34345 38845 34379 38879
rect 34462 38845 34496 38879
rect 34621 38845 34655 38879
rect 41797 38845 41831 38879
rect 42625 38845 42659 38879
rect 42809 38845 42843 38879
rect 50629 38845 50663 38879
rect 34069 38777 34103 38811
rect 20637 38709 20671 38743
rect 32505 38709 32539 38743
rect 36001 38709 36035 38743
rect 36553 38709 36587 38743
rect 23673 38505 23707 38539
rect 27721 38505 27755 38539
rect 32781 38505 32815 38539
rect 36921 38505 36955 38539
rect 41613 38505 41647 38539
rect 44281 38437 44315 38471
rect 37381 38369 37415 38403
rect 45845 38369 45879 38403
rect 46029 38369 46063 38403
rect 19809 38301 19843 38335
rect 20913 38301 20947 38335
rect 23581 38301 23615 38335
rect 24409 38301 24443 38335
rect 27905 38301 27939 38335
rect 29837 38301 29871 38335
rect 30849 38301 30883 38335
rect 30941 38301 30975 38335
rect 31401 38301 31435 38335
rect 34989 38301 35023 38335
rect 35081 38301 35115 38335
rect 35541 38301 35575 38335
rect 35808 38301 35842 38335
rect 37657 38301 37691 38335
rect 40417 38301 40451 38335
rect 42165 38301 42199 38335
rect 42441 38301 42475 38335
rect 42901 38301 42935 38335
rect 43168 38301 43202 38335
rect 50169 38301 50203 38335
rect 21180 38233 21214 38267
rect 24676 38233 24710 38267
rect 31668 38233 31702 38267
rect 33793 38233 33827 38267
rect 33977 38233 34011 38267
rect 40601 38233 40635 38267
rect 41521 38233 41555 38267
rect 47685 38233 47719 38267
rect 19901 38165 19935 38199
rect 22293 38165 22327 38199
rect 25789 38165 25823 38199
rect 29653 38165 29687 38199
rect 50261 38165 50295 38199
rect 25329 37961 25363 37995
rect 32137 37961 32171 37995
rect 19625 37893 19659 37927
rect 27169 37893 27203 37927
rect 27385 37893 27419 37927
rect 29644 37893 29678 37927
rect 37749 37893 37783 37927
rect 38761 37893 38795 37927
rect 40110 37893 40144 37927
rect 44373 37893 44407 37927
rect 50077 37893 50111 37927
rect 19441 37825 19475 37859
rect 23305 37825 23339 37859
rect 25329 37825 25363 37859
rect 26065 37825 26099 37859
rect 29377 37825 29411 37859
rect 32321 37825 32355 37859
rect 32873 37825 32907 37859
rect 35541 37825 35575 37859
rect 37565 37825 37599 37859
rect 39017 37825 39051 37859
rect 39129 37825 39163 37859
rect 39221 37828 39255 37862
rect 39405 37825 39439 37859
rect 39865 37825 39899 37859
rect 42441 37825 42475 37859
rect 42717 37825 42751 37859
rect 45017 37825 45051 37859
rect 19901 37757 19935 37791
rect 24225 37757 24259 37791
rect 33149 37757 33183 37791
rect 35725 37757 35759 37791
rect 47593 37757 47627 37791
rect 47777 37757 47811 37791
rect 48053 37757 48087 37791
rect 49893 37757 49927 37791
rect 51733 37757 51767 37791
rect 37933 37689 37967 37723
rect 41245 37689 41279 37723
rect 25881 37621 25915 37655
rect 27353 37621 27387 37655
rect 27537 37621 27571 37655
rect 30757 37621 30791 37655
rect 44465 37621 44499 37655
rect 45201 37621 45235 37655
rect 29009 37417 29043 37451
rect 38761 37417 38795 37451
rect 47317 37417 47351 37451
rect 26709 37349 26743 37383
rect 27813 37349 27847 37383
rect 22477 37281 22511 37315
rect 24501 37281 24535 37315
rect 25329 37281 25363 37315
rect 27169 37281 27203 37315
rect 28206 37281 28240 37315
rect 29745 37281 29779 37315
rect 35449 37281 35483 37315
rect 39129 37281 39163 37315
rect 41153 37281 41187 37315
rect 41613 37281 41647 37315
rect 22017 37213 22051 37247
rect 24685 37213 24719 37247
rect 27353 37213 27387 37247
rect 28089 37213 28123 37247
rect 28365 37213 28399 37247
rect 30021 37213 30055 37247
rect 32781 37213 32815 37247
rect 34897 37213 34931 37247
rect 35725 37213 35759 37247
rect 36737 37213 36771 37247
rect 38945 37213 38979 37247
rect 39037 37213 39071 37247
rect 39221 37213 39255 37247
rect 40969 37213 41003 37247
rect 41889 37213 41923 37247
rect 42993 37213 43027 37247
rect 44097 37213 44131 37247
rect 45201 37213 45235 37247
rect 47225 37213 47259 37247
rect 22201 37145 22235 37179
rect 25596 37145 25630 37179
rect 33048 37145 33082 37179
rect 43177 37145 43211 37179
rect 44281 37145 44315 37179
rect 45446 37145 45480 37179
rect 24869 37077 24903 37111
rect 34161 37077 34195 37111
rect 34713 37077 34747 37111
rect 36921 37077 36955 37111
rect 46581 37077 46615 37111
rect 22753 36873 22787 36907
rect 24685 36873 24719 36907
rect 30037 36873 30071 36907
rect 30205 36873 30239 36907
rect 39405 36873 39439 36907
rect 44833 36873 44867 36907
rect 29837 36805 29871 36839
rect 36185 36805 36219 36839
rect 36385 36805 36419 36839
rect 37565 36805 37599 36839
rect 37749 36805 37783 36839
rect 40693 36805 40727 36839
rect 43913 36805 43947 36839
rect 2513 36737 2547 36771
rect 22661 36737 22695 36771
rect 23397 36737 23431 36771
rect 24869 36737 24903 36771
rect 25881 36737 25915 36771
rect 27261 36737 27295 36771
rect 30757 36737 30791 36771
rect 32597 36737 32631 36771
rect 32873 36737 32907 36771
rect 33885 36737 33919 36771
rect 34069 36737 34103 36771
rect 37381 36737 37415 36771
rect 38209 36737 38243 36771
rect 38393 36737 38427 36771
rect 39037 36737 39071 36771
rect 39221 36737 39255 36771
rect 41613 36737 41647 36771
rect 41705 36737 41739 36771
rect 43177 36737 43211 36771
rect 43269 36737 43303 36771
rect 44097 36737 44131 36771
rect 45089 36737 45123 36771
rect 45182 36740 45216 36774
rect 45282 36737 45316 36771
rect 45477 36737 45511 36771
rect 46213 36737 46247 36771
rect 46305 36737 46339 36771
rect 46397 36737 46431 36771
rect 46581 36737 46615 36771
rect 25605 36669 25639 36703
rect 27537 36669 27571 36703
rect 28549 36669 28583 36703
rect 28825 36669 28859 36703
rect 31033 36669 31067 36703
rect 34805 36669 34839 36703
rect 34922 36669 34956 36703
rect 35081 36669 35115 36703
rect 35725 36669 35759 36703
rect 38577 36669 38611 36703
rect 41521 36669 41555 36703
rect 41797 36669 41831 36703
rect 43085 36669 43119 36703
rect 43361 36669 43395 36703
rect 34529 36601 34563 36635
rect 44281 36601 44315 36635
rect 2605 36533 2639 36567
rect 23673 36533 23707 36567
rect 30021 36533 30055 36567
rect 36369 36533 36403 36567
rect 36553 36533 36587 36567
rect 40785 36533 40819 36567
rect 41337 36533 41371 36567
rect 42901 36533 42935 36567
rect 45937 36533 45971 36567
rect 26617 36329 26651 36363
rect 32321 36329 32355 36363
rect 33333 36329 33367 36363
rect 33517 36329 33551 36363
rect 37381 36329 37415 36363
rect 39313 36329 39347 36363
rect 47869 36329 47903 36363
rect 23673 36261 23707 36295
rect 1593 36193 1627 36227
rect 2789 36193 2823 36227
rect 24409 36193 24443 36227
rect 36001 36193 36035 36227
rect 40141 36193 40175 36227
rect 43361 36193 43395 36227
rect 1409 36125 1443 36159
rect 22293 36125 22327 36159
rect 24593 36125 24627 36159
rect 25237 36125 25271 36159
rect 26801 36125 26835 36159
rect 28549 36125 28583 36159
rect 29745 36125 29779 36159
rect 30297 36125 30331 36159
rect 30481 36125 30515 36159
rect 30941 36125 30975 36159
rect 37933 36125 37967 36159
rect 39865 36125 39899 36159
rect 41521 36125 41555 36159
rect 41797 36125 41831 36159
rect 43545 36125 43579 36159
rect 46489 36125 46523 36159
rect 46745 36125 46779 36159
rect 67925 36125 67959 36159
rect 22560 36057 22594 36091
rect 31208 36057 31242 36091
rect 33149 36057 33183 36091
rect 36268 36057 36302 36091
rect 38200 36057 38234 36091
rect 24777 35989 24811 36023
rect 25329 35989 25363 36023
rect 28733 35989 28767 36023
rect 29561 35989 29595 36023
rect 33349 35989 33383 36023
rect 43729 35989 43763 36023
rect 19717 35785 19751 35819
rect 23213 35785 23247 35819
rect 36369 35785 36403 35819
rect 38393 35785 38427 35819
rect 20085 35717 20119 35751
rect 28908 35717 28942 35751
rect 42441 35717 42475 35751
rect 42809 35717 42843 35751
rect 46949 35717 46983 35751
rect 48145 35717 48179 35751
rect 2145 35649 2179 35683
rect 19165 35649 19199 35683
rect 19533 35649 19567 35683
rect 20729 35649 20763 35683
rect 21005 35649 21039 35683
rect 21833 35649 21867 35683
rect 22477 35649 22511 35683
rect 22661 35649 22695 35683
rect 23029 35649 23063 35683
rect 24225 35649 24259 35683
rect 24492 35649 24526 35683
rect 27169 35649 27203 35683
rect 28641 35649 28675 35683
rect 30481 35649 30515 35683
rect 31309 35649 31343 35683
rect 31401 35649 31435 35683
rect 32413 35649 32447 35683
rect 33333 35649 33367 35683
rect 35173 35649 35207 35683
rect 35633 35649 35667 35683
rect 36553 35649 36587 35683
rect 38209 35649 38243 35683
rect 39221 35649 39255 35683
rect 39313 35649 39347 35683
rect 40776 35649 40810 35683
rect 42625 35649 42659 35683
rect 43720 35649 43754 35683
rect 46857 35649 46891 35683
rect 47961 35649 47995 35683
rect 65809 35649 65843 35683
rect 19073 35581 19107 35615
rect 20913 35581 20947 35615
rect 40509 35581 40543 35615
rect 43453 35581 43487 35615
rect 49617 35581 49651 35615
rect 65993 35581 66027 35615
rect 67557 35581 67591 35615
rect 21189 35513 21223 35547
rect 30665 35513 30699 35547
rect 35633 35513 35667 35547
rect 41889 35513 41923 35547
rect 44833 35513 44867 35547
rect 19533 35445 19567 35479
rect 20453 35445 20487 35479
rect 21005 35445 21039 35479
rect 25605 35445 25639 35479
rect 26985 35445 27019 35479
rect 30021 35445 30055 35479
rect 31585 35445 31619 35479
rect 32597 35445 32631 35479
rect 33149 35445 33183 35479
rect 34989 35445 35023 35479
rect 39497 35445 39531 35479
rect 20177 35241 20211 35275
rect 20637 35241 20671 35275
rect 22293 35241 22327 35275
rect 23029 35241 23063 35275
rect 29745 35241 29779 35275
rect 29929 35241 29963 35275
rect 31309 35241 31343 35275
rect 36553 35241 36587 35275
rect 38945 35241 38979 35275
rect 43637 35241 43671 35275
rect 67557 35241 67591 35275
rect 21005 35173 21039 35207
rect 26709 35173 26743 35207
rect 27813 35173 27847 35207
rect 35357 35173 35391 35207
rect 45661 35173 45695 35207
rect 20637 35105 20671 35139
rect 24501 35105 24535 35139
rect 27169 35105 27203 35139
rect 27353 35105 27387 35139
rect 28206 35105 28240 35139
rect 32597 35105 32631 35139
rect 34897 35105 34931 35139
rect 35750 35105 35784 35139
rect 35909 35105 35943 35139
rect 40141 35105 40175 35139
rect 40417 35105 40451 35139
rect 41521 35105 41555 35139
rect 42809 35105 42843 35139
rect 49249 35105 49283 35139
rect 20821 35037 20855 35071
rect 22385 35037 22419 35071
rect 23213 35037 23247 35071
rect 24685 35037 24719 35071
rect 25329 35037 25363 35071
rect 25596 35037 25630 35071
rect 28089 35037 28123 35071
rect 28365 35037 28399 35071
rect 29009 35037 29043 35071
rect 30573 35037 30607 35071
rect 31493 35037 31527 35071
rect 32864 35037 32898 35071
rect 34713 35037 34747 35071
rect 35633 35037 35667 35071
rect 38485 35037 38519 35071
rect 39129 35037 39163 35071
rect 41797 35037 41831 35071
rect 42993 35037 43027 35071
rect 43637 35037 43671 35071
rect 45477 35037 45511 35071
rect 47501 35037 47535 35071
rect 67465 35037 67499 35071
rect 20545 34969 20579 35003
rect 29561 34969 29595 35003
rect 37197 34969 37231 35003
rect 37381 34969 37415 35003
rect 47685 34969 47719 35003
rect 24869 34901 24903 34935
rect 29761 34901 29795 34935
rect 30573 34901 30607 34935
rect 33977 34901 34011 34935
rect 37565 34901 37599 34935
rect 38301 34901 38335 34935
rect 43177 34901 43211 34935
rect 24685 34697 24719 34731
rect 25973 34697 26007 34731
rect 27445 34697 27479 34731
rect 31585 34697 31619 34731
rect 32137 34697 32171 34731
rect 33425 34697 33459 34731
rect 36737 34697 36771 34731
rect 38945 34697 38979 34731
rect 40969 34697 41003 34731
rect 41613 34697 41647 34731
rect 44005 34697 44039 34731
rect 46857 34697 46891 34731
rect 47685 34697 47719 34731
rect 27077 34629 27111 34663
rect 27293 34629 27327 34663
rect 30472 34629 30506 34663
rect 33057 34629 33091 34663
rect 33257 34629 33291 34663
rect 37749 34629 37783 34663
rect 1685 34561 1719 34595
rect 23121 34561 23155 34595
rect 24869 34561 24903 34595
rect 25973 34561 26007 34595
rect 30205 34561 30239 34595
rect 32321 34561 32355 34595
rect 35357 34561 35391 34595
rect 35613 34561 35647 34595
rect 39221 34561 39255 34595
rect 39313 34561 39347 34595
rect 40969 34561 41003 34595
rect 41797 34561 41831 34595
rect 44189 34561 44223 34595
rect 45477 34561 45511 34595
rect 45744 34561 45778 34595
rect 47593 34561 47627 34595
rect 67281 34561 67315 34595
rect 1409 34493 1443 34527
rect 39129 34493 39163 34527
rect 39405 34493 39439 34527
rect 22937 34357 22971 34391
rect 27261 34357 27295 34391
rect 33241 34357 33275 34391
rect 37841 34357 37875 34391
rect 67373 34357 67407 34391
rect 23857 34153 23891 34187
rect 28549 34153 28583 34187
rect 30481 34153 30515 34187
rect 31493 34153 31527 34187
rect 35817 34153 35851 34187
rect 36001 34153 36035 34187
rect 45109 34153 45143 34187
rect 31125 34017 31159 34051
rect 40417 34017 40451 34051
rect 42717 34017 42751 34051
rect 42901 34017 42935 34051
rect 22477 33949 22511 33983
rect 22744 33949 22778 33983
rect 24593 33949 24627 33983
rect 25329 33949 25363 33983
rect 28365 33949 28399 33983
rect 29561 33949 29595 33983
rect 30297 33949 30331 33983
rect 31309 33949 31343 33983
rect 37197 33949 37231 33983
rect 37381 33949 37415 33983
rect 37841 33949 37875 33983
rect 38108 33949 38142 33983
rect 42809 33949 42843 33983
rect 42993 33949 43027 33983
rect 43913 33949 43947 33983
rect 45385 33949 45419 33983
rect 45477 33949 45511 33983
rect 45569 33949 45603 33983
rect 45753 33949 45787 33983
rect 35633 33881 35667 33915
rect 40662 33881 40696 33915
rect 24593 33813 24627 33847
rect 25145 33813 25179 33847
rect 29745 33813 29779 33847
rect 35833 33813 35867 33847
rect 39221 33813 39255 33847
rect 41797 33813 41831 33847
rect 42533 33813 42567 33847
rect 43729 33813 43763 33847
rect 22569 33609 22603 33643
rect 23489 33609 23523 33643
rect 38485 33609 38519 33643
rect 40049 33609 40083 33643
rect 43177 33609 43211 33643
rect 45017 33609 45051 33643
rect 24676 33541 24710 33575
rect 32965 33541 32999 33575
rect 33181 33541 33215 33575
rect 38117 33541 38151 33575
rect 39313 33541 39347 33575
rect 43882 33541 43916 33575
rect 22385 33473 22419 33507
rect 23213 33473 23247 33507
rect 23305 33473 23339 33507
rect 24409 33473 24443 33507
rect 27537 33473 27571 33507
rect 28549 33473 28583 33507
rect 29653 33473 29687 33507
rect 30481 33473 30515 33507
rect 35633 33473 35667 33507
rect 38301 33473 38335 33507
rect 39037 33473 39071 33507
rect 39129 33473 39163 33507
rect 40325 33473 40359 33507
rect 40417 33473 40451 33507
rect 40509 33473 40543 33507
rect 40693 33473 40727 33507
rect 42901 33473 42935 33507
rect 42993 33473 43027 33507
rect 46857 33473 46891 33507
rect 27353 33405 27387 33439
rect 27997 33405 28031 33439
rect 28273 33405 28307 33439
rect 28390 33405 28424 33439
rect 35357 33405 35391 33439
rect 43637 33405 43671 33439
rect 29193 33337 29227 33371
rect 25789 33269 25823 33303
rect 29837 33269 29871 33303
rect 30573 33269 30607 33303
rect 33149 33269 33183 33303
rect 33333 33269 33367 33303
rect 46949 33269 46983 33303
rect 67649 33269 67683 33303
rect 24961 33065 24995 33099
rect 27629 33065 27663 33099
rect 28273 33065 28307 33099
rect 33793 33065 33827 33099
rect 34897 33065 34931 33099
rect 42993 33065 43027 33099
rect 43637 33065 43671 33099
rect 36921 32997 36955 33031
rect 46949 32929 46983 32963
rect 66269 32929 66303 32963
rect 23029 32861 23063 32895
rect 26249 32861 26283 32895
rect 29745 32861 29779 32895
rect 31125 32861 31159 32895
rect 32413 32861 32447 32895
rect 35541 32861 35575 32895
rect 37381 32861 37415 32895
rect 37565 32861 37599 32895
rect 38669 32861 38703 32895
rect 42625 32861 42659 32895
rect 42809 32861 42843 32895
rect 43453 32861 43487 32895
rect 44281 32861 44315 32895
rect 46765 32861 46799 32895
rect 24869 32793 24903 32827
rect 26516 32793 26550 32827
rect 28089 32793 28123 32827
rect 28305 32793 28339 32827
rect 32680 32793 32714 32827
rect 34713 32793 34747 32827
rect 35808 32793 35842 32827
rect 48605 32793 48639 32827
rect 66453 32793 66487 32827
rect 68109 32793 68143 32827
rect 22845 32725 22879 32759
rect 28457 32725 28491 32759
rect 29561 32725 29595 32759
rect 30941 32725 30975 32759
rect 34913 32725 34947 32759
rect 35081 32725 35115 32759
rect 37749 32725 37783 32759
rect 38761 32725 38795 32759
rect 44373 32725 44407 32759
rect 25697 32521 25731 32555
rect 26341 32521 26375 32555
rect 26985 32521 27019 32555
rect 30113 32521 30147 32555
rect 31401 32521 31435 32555
rect 32413 32521 32447 32555
rect 36461 32521 36495 32555
rect 44097 32521 44131 32555
rect 67557 32521 67591 32555
rect 22652 32453 22686 32487
rect 29000 32453 29034 32487
rect 35265 32453 35299 32487
rect 37289 32453 37323 32487
rect 37473 32453 37507 32487
rect 42901 32453 42935 32487
rect 25421 32385 25455 32419
rect 25513 32385 25547 32419
rect 26157 32385 26191 32419
rect 27169 32385 27203 32419
rect 31217 32385 31251 32419
rect 32321 32385 32355 32419
rect 33425 32385 33459 32419
rect 35817 32385 35851 32419
rect 36645 32385 36679 32419
rect 38393 32385 38427 32419
rect 38577 32385 38611 32419
rect 39313 32385 39347 32419
rect 39580 32385 39614 32419
rect 41245 32385 41279 32419
rect 42717 32385 42751 32419
rect 44373 32385 44407 32419
rect 44462 32385 44496 32419
rect 44557 32385 44591 32419
rect 44741 32385 44775 32419
rect 45468 32385 45502 32419
rect 67465 32385 67499 32419
rect 22385 32317 22419 32351
rect 28733 32317 28767 32351
rect 31033 32317 31067 32351
rect 33609 32317 33643 32351
rect 34345 32317 34379 32351
rect 34462 32317 34496 32351
rect 34621 32317 34655 32351
rect 38301 32317 38335 32351
rect 38485 32317 38519 32351
rect 45201 32317 45235 32351
rect 23765 32249 23799 32283
rect 34069 32249 34103 32283
rect 37657 32249 37691 32283
rect 35909 32181 35943 32215
rect 38117 32181 38151 32215
rect 40693 32181 40727 32215
rect 41429 32181 41463 32215
rect 43085 32181 43119 32215
rect 46581 32181 46615 32215
rect 22477 31977 22511 32011
rect 23397 31977 23431 32011
rect 28825 31977 28859 32011
rect 29745 31977 29779 32011
rect 29929 31977 29963 32011
rect 32873 31977 32907 32011
rect 35633 31977 35667 32011
rect 39221 31977 39255 32011
rect 43177 31977 43211 32011
rect 31953 31909 31987 31943
rect 37289 31909 37323 31943
rect 42717 31909 42751 31943
rect 23029 31841 23063 31875
rect 24777 31841 24811 31875
rect 30573 31841 30607 31875
rect 39865 31841 39899 31875
rect 41337 31841 41371 31875
rect 43453 31841 43487 31875
rect 43545 31841 43579 31875
rect 43637 31841 43671 31875
rect 1869 31773 1903 31807
rect 22477 31773 22511 31807
rect 23213 31773 23247 31807
rect 24501 31773 24535 31807
rect 25973 31773 26007 31807
rect 26709 31773 26743 31807
rect 28641 31773 28675 31807
rect 30840 31773 30874 31807
rect 33057 31773 33091 31807
rect 35633 31773 35667 31807
rect 36921 31773 36955 31807
rect 37105 31773 37139 31807
rect 38853 31773 38887 31807
rect 39037 31773 39071 31807
rect 40049 31773 40083 31807
rect 43361 31773 43395 31807
rect 67925 31773 67959 31807
rect 29561 31705 29595 31739
rect 29761 31705 29795 31739
rect 41604 31705 41638 31739
rect 25973 31637 26007 31671
rect 26525 31637 26559 31671
rect 40233 31637 40267 31671
rect 23213 31433 23247 31467
rect 27353 31433 27387 31467
rect 28013 31433 28047 31467
rect 39681 31433 39715 31467
rect 41705 31433 41739 31467
rect 25320 31365 25354 31399
rect 26985 31365 27019 31399
rect 27201 31365 27235 31399
rect 27813 31365 27847 31399
rect 35357 31365 35391 31399
rect 35557 31365 35591 31399
rect 38853 31365 38887 31399
rect 1685 31297 1719 31331
rect 23029 31297 23063 31331
rect 25053 31297 25087 31331
rect 31585 31297 31619 31331
rect 32413 31297 32447 31331
rect 33416 31297 33450 31331
rect 36185 31297 36219 31331
rect 37749 31297 37783 31331
rect 39037 31297 39071 31331
rect 39865 31297 39899 31331
rect 41889 31297 41923 31331
rect 42533 31297 42567 31331
rect 42625 31297 42659 31331
rect 43729 31297 43763 31331
rect 44649 31297 44683 31331
rect 65809 31297 65843 31331
rect 1869 31229 1903 31263
rect 2789 31229 2823 31263
rect 32689 31229 32723 31263
rect 33149 31229 33183 31263
rect 42809 31229 42843 31263
rect 65993 31229 66027 31263
rect 67557 31229 67591 31263
rect 26433 31093 26467 31127
rect 27169 31093 27203 31127
rect 27997 31093 28031 31127
rect 28181 31093 28215 31127
rect 31401 31093 31435 31127
rect 34529 31093 34563 31127
rect 35541 31093 35575 31127
rect 35725 31093 35759 31127
rect 36185 31093 36219 31127
rect 37565 31093 37599 31127
rect 39221 31093 39255 31127
rect 43913 31093 43947 31127
rect 44465 31093 44499 31127
rect 2053 30889 2087 30923
rect 33425 30889 33459 30923
rect 34713 30889 34747 30923
rect 44189 30889 44223 30923
rect 67649 30889 67683 30923
rect 33609 30821 33643 30855
rect 37565 30753 37599 30787
rect 1961 30685 1995 30719
rect 22477 30685 22511 30719
rect 23213 30685 23247 30719
rect 24593 30685 24627 30719
rect 28549 30685 28583 30719
rect 29561 30685 29595 30719
rect 31125 30685 31159 30719
rect 31392 30685 31426 30719
rect 34897 30685 34931 30719
rect 35541 30685 35575 30719
rect 40417 30685 40451 30719
rect 40601 30685 40635 30719
rect 41245 30685 41279 30719
rect 42993 30685 43027 30719
rect 43913 30685 43947 30719
rect 44005 30685 44039 30719
rect 67557 30685 67591 30719
rect 23397 30617 23431 30651
rect 33241 30617 33275 30651
rect 33441 30617 33475 30651
rect 35786 30617 35820 30651
rect 37832 30617 37866 30651
rect 43177 30617 43211 30651
rect 22293 30549 22327 30583
rect 24409 30549 24443 30583
rect 28365 30549 28399 30583
rect 29653 30549 29687 30583
rect 32505 30549 32539 30583
rect 36921 30549 36955 30583
rect 38945 30549 38979 30583
rect 40785 30549 40819 30583
rect 41429 30549 41463 30583
rect 43361 30549 43395 30583
rect 23029 30345 23063 30379
rect 31125 30345 31159 30379
rect 32965 30345 32999 30379
rect 38209 30345 38243 30379
rect 41889 30345 41923 30379
rect 45477 30345 45511 30379
rect 23756 30277 23790 30311
rect 28794 30277 28828 30311
rect 32597 30277 32631 30311
rect 32813 30277 32847 30311
rect 36553 30277 36587 30311
rect 37473 30277 37507 30311
rect 44364 30277 44398 30311
rect 22017 30209 22051 30243
rect 22845 30209 22879 30243
rect 23489 30209 23523 30243
rect 28549 30209 28583 30243
rect 31125 30209 31159 30243
rect 33517 30209 33551 30243
rect 33701 30209 33735 30243
rect 35357 30209 35391 30243
rect 36369 30209 36403 30243
rect 37289 30209 37323 30243
rect 38393 30209 38427 30243
rect 39129 30209 39163 30243
rect 39313 30209 39347 30243
rect 40509 30209 40543 30243
rect 40765 30209 40799 30243
rect 42993 30209 43027 30243
rect 43177 30209 43211 30243
rect 44097 30209 44131 30243
rect 1869 30141 1903 30175
rect 2053 30141 2087 30175
rect 2881 30141 2915 30175
rect 22661 30141 22695 30175
rect 34437 30141 34471 30175
rect 34554 30141 34588 30175
rect 34713 30141 34747 30175
rect 37657 30141 37691 30175
rect 39221 30141 39255 30175
rect 39405 30141 39439 30175
rect 43085 30141 43119 30175
rect 43269 30141 43303 30175
rect 34161 30073 34195 30107
rect 36737 30073 36771 30107
rect 21925 30005 21959 30039
rect 24869 30005 24903 30039
rect 29929 30005 29963 30039
rect 32781 30005 32815 30039
rect 38945 30005 38979 30039
rect 42809 30005 42843 30039
rect 2053 29801 2087 29835
rect 2789 29801 2823 29835
rect 23213 29801 23247 29835
rect 24777 29801 24811 29835
rect 28273 29801 28307 29835
rect 35357 29801 35391 29835
rect 39129 29801 39163 29835
rect 27077 29733 27111 29767
rect 31125 29733 31159 29767
rect 21833 29665 21867 29699
rect 24409 29665 24443 29699
rect 26433 29665 26467 29699
rect 27470 29665 27504 29699
rect 27629 29665 27663 29699
rect 31585 29665 31619 29699
rect 37197 29665 37231 29699
rect 40969 29665 41003 29699
rect 41061 29665 41095 29699
rect 2697 29597 2731 29631
rect 22100 29597 22134 29631
rect 24593 29597 24627 29631
rect 25421 29597 25455 29631
rect 26617 29597 26651 29631
rect 27353 29597 27387 29631
rect 29745 29597 29779 29631
rect 31769 29597 31803 29631
rect 35541 29597 35575 29631
rect 37013 29597 37047 29631
rect 38853 29597 38887 29631
rect 38945 29597 38979 29631
rect 39865 29597 39899 29631
rect 40049 29597 40083 29631
rect 40233 29597 40267 29631
rect 40877 29597 40911 29631
rect 41153 29597 41187 29631
rect 45017 29597 45051 29631
rect 30012 29529 30046 29563
rect 36829 29529 36863 29563
rect 25237 29461 25271 29495
rect 31953 29461 31987 29495
rect 40693 29461 40727 29495
rect 45109 29461 45143 29495
rect 29009 29257 29043 29291
rect 29653 29257 29687 29291
rect 30297 29257 30331 29291
rect 33977 29257 34011 29291
rect 35281 29257 35315 29291
rect 35449 29257 35483 29291
rect 40601 29257 40635 29291
rect 24952 29189 24986 29223
rect 35081 29189 35115 29223
rect 44281 29189 44315 29223
rect 27169 29121 27203 29155
rect 28089 29121 28123 29155
rect 29653 29121 29687 29155
rect 30481 29121 30515 29155
rect 32137 29121 32171 29155
rect 32321 29121 32355 29155
rect 36093 29121 36127 29155
rect 38209 29121 38243 29155
rect 38301 29121 38335 29155
rect 38393 29121 38427 29155
rect 38577 29121 38611 29155
rect 39313 29121 39347 29155
rect 39405 29121 39439 29155
rect 39497 29121 39531 29155
rect 39681 29121 39715 29155
rect 40785 29121 40819 29155
rect 43085 29121 43119 29155
rect 43177 29121 43211 29155
rect 43269 29121 43303 29155
rect 43453 29121 43487 29155
rect 24685 29053 24719 29087
rect 27353 29053 27387 29087
rect 28206 29053 28240 29087
rect 28365 29053 28399 29087
rect 33057 29053 33091 29087
rect 33174 29053 33208 29087
rect 33333 29053 33367 29087
rect 44097 29053 44131 29087
rect 45937 29053 45971 29087
rect 27813 28985 27847 29019
rect 32781 28985 32815 29019
rect 26065 28917 26099 28951
rect 35265 28917 35299 28951
rect 35909 28917 35943 28951
rect 37933 28917 37967 28951
rect 39037 28917 39071 28951
rect 42809 28917 42843 28951
rect 24777 28713 24811 28747
rect 25697 28713 25731 28747
rect 36553 28713 36587 28747
rect 44189 28713 44223 28747
rect 25329 28577 25363 28611
rect 31217 28577 31251 28611
rect 40969 28577 41003 28611
rect 24777 28509 24811 28543
rect 25513 28509 25547 28543
rect 26341 28509 26375 28543
rect 29745 28509 29779 28543
rect 31401 28509 31435 28543
rect 35173 28509 35207 28543
rect 35440 28509 35474 28543
rect 37013 28509 37047 28543
rect 42809 28509 42843 28543
rect 43065 28509 43099 28543
rect 37280 28441 37314 28475
rect 41214 28441 41248 28475
rect 26341 28373 26375 28407
rect 29929 28373 29963 28407
rect 31585 28373 31619 28407
rect 38393 28373 38427 28407
rect 42349 28373 42383 28407
rect 35541 28169 35575 28203
rect 40877 28169 40911 28203
rect 27997 28101 28031 28135
rect 28213 28101 28247 28135
rect 28825 28101 28859 28135
rect 29041 28101 29075 28135
rect 23029 28033 23063 28067
rect 25697 28033 25731 28067
rect 25881 28033 25915 28067
rect 27169 28033 27203 28067
rect 30205 28033 30239 28067
rect 30472 28033 30506 28067
rect 33425 28033 33459 28067
rect 35357 28033 35391 28067
rect 38853 28033 38887 28067
rect 39120 28033 39154 28067
rect 41153 28033 41187 28067
rect 41245 28033 41279 28067
rect 41337 28033 41371 28067
rect 41521 28033 41555 28067
rect 23213 27965 23247 27999
rect 23489 27965 23523 27999
rect 25513 27965 25547 27999
rect 34069 27965 34103 27999
rect 34345 27965 34379 27999
rect 31585 27897 31619 27931
rect 26985 27829 27019 27863
rect 28181 27829 28215 27863
rect 28365 27829 28399 27863
rect 29009 27829 29043 27863
rect 29193 27829 29227 27863
rect 33241 27829 33275 27863
rect 40233 27829 40267 27863
rect 23213 27625 23247 27659
rect 28365 27625 28399 27659
rect 31217 27625 31251 27659
rect 34069 27557 34103 27591
rect 35081 27557 35115 27591
rect 26157 27489 26191 27523
rect 34713 27489 34747 27523
rect 37197 27489 37231 27523
rect 38577 27489 38611 27523
rect 23121 27421 23155 27455
rect 24409 27421 24443 27455
rect 26985 27421 27019 27455
rect 29009 27421 29043 27455
rect 29745 27421 29779 27455
rect 30481 27421 30515 27455
rect 31401 27421 31435 27455
rect 32689 27421 32723 27455
rect 32956 27421 32990 27455
rect 34897 27421 34931 27455
rect 40877 27421 40911 27455
rect 24593 27353 24627 27387
rect 27252 27353 27286 27387
rect 37381 27353 37415 27387
rect 28825 27285 28859 27319
rect 29745 27285 29779 27319
rect 30665 27285 30699 27319
rect 40969 27285 41003 27319
rect 24501 27081 24535 27115
rect 26433 27081 26467 27115
rect 27629 27081 27663 27115
rect 30021 27081 30055 27115
rect 32689 27081 32723 27115
rect 36001 27081 36035 27115
rect 37381 27081 37415 27115
rect 25320 27013 25354 27047
rect 24409 26945 24443 26979
rect 25053 26945 25087 26979
rect 27537 26945 27571 26979
rect 28641 26945 28675 26979
rect 28908 26945 28942 26979
rect 32505 26945 32539 26979
rect 33977 26945 34011 26979
rect 34621 26945 34655 26979
rect 34888 26945 34922 26979
rect 37289 26945 37323 26979
rect 40049 26945 40083 26979
rect 33793 26877 33827 26911
rect 40233 26877 40267 26911
rect 40509 26877 40543 26911
rect 34161 26741 34195 26775
rect 27537 26537 27571 26571
rect 34713 26537 34747 26571
rect 35449 26537 35483 26571
rect 40325 26537 40359 26571
rect 32505 26469 32539 26503
rect 32965 26401 32999 26435
rect 41337 26401 41371 26435
rect 41521 26401 41555 26435
rect 1961 26333 1995 26367
rect 27721 26333 27755 26367
rect 31125 26333 31159 26367
rect 33149 26333 33183 26367
rect 34713 26333 34747 26367
rect 35633 26333 35667 26367
rect 40233 26333 40267 26367
rect 31392 26265 31426 26299
rect 43177 26265 43211 26299
rect 33333 26197 33367 26231
rect 31125 25993 31159 26027
rect 32137 25993 32171 26027
rect 35081 25993 35115 26027
rect 1685 25857 1719 25891
rect 31125 25857 31159 25891
rect 32321 25857 32355 25891
rect 33968 25857 34002 25891
rect 1869 25789 1903 25823
rect 2789 25789 2823 25823
rect 33701 25789 33735 25823
rect 2329 25449 2363 25483
rect 33793 25449 33827 25483
rect 32505 25313 32539 25347
rect 2237 25245 2271 25279
rect 32689 25245 32723 25279
rect 33793 25245 33827 25279
rect 34805 25245 34839 25279
rect 34897 25245 34931 25279
rect 32873 25109 32907 25143
rect 35081 25109 35115 25143
rect 34069 24905 34103 24939
rect 1869 24769 1903 24803
rect 2605 24769 2639 24803
rect 31401 24769 31435 24803
rect 32393 24769 32427 24803
rect 34253 24769 34287 24803
rect 2053 24701 2087 24735
rect 31493 24701 31527 24735
rect 32137 24701 32171 24735
rect 2697 24565 2731 24599
rect 3433 24565 3467 24599
rect 33517 24565 33551 24599
rect 32229 24361 32263 24395
rect 1409 24225 1443 24259
rect 1593 24225 1627 24259
rect 2789 24225 2823 24259
rect 32413 24157 32447 24191
rect 67649 23477 67683 23511
rect 66269 23137 66303 23171
rect 68109 23137 68143 23171
rect 66453 23001 66487 23035
rect 67281 22729 67315 22763
rect 67189 22593 67223 22627
rect 1777 22525 1811 22559
rect 1961 22525 1995 22559
rect 2789 22525 2823 22559
rect 2053 22185 2087 22219
rect 2605 22185 2639 22219
rect 67925 22117 67959 22151
rect 2513 21981 2547 22015
rect 65993 21573 66027 21607
rect 1869 21505 1903 21539
rect 65809 21437 65843 21471
rect 67557 21437 67591 21471
rect 1961 21301 1995 21335
rect 67833 18717 67867 18751
rect 68017 18581 68051 18615
rect 27721 18309 27755 18343
rect 26985 18241 27019 18275
rect 27353 18173 27387 18207
rect 27261 18105 27295 18139
rect 27150 18037 27184 18071
rect 67925 17629 67959 17663
rect 65993 17221 66027 17255
rect 65809 17153 65843 17187
rect 67557 17085 67591 17119
rect 67557 16541 67591 16575
rect 67649 16405 67683 16439
rect 2053 15997 2087 16031
rect 2237 15997 2271 16031
rect 2973 15997 3007 16031
rect 2329 15657 2363 15691
rect 2881 15657 2915 15691
rect 2789 15453 2823 15487
rect 67557 15453 67591 15487
rect 67649 15317 67683 15351
rect 65993 15045 66027 15079
rect 65809 14909 65843 14943
rect 67557 14909 67591 14943
rect 67925 14569 67959 14603
rect 1777 13277 1811 13311
rect 67833 13277 67867 13311
rect 68017 13141 68051 13175
rect 1593 12801 1627 12835
rect 32137 12801 32171 12835
rect 33149 12801 33183 12835
rect 1777 12733 1811 12767
rect 2789 12733 2823 12767
rect 32284 12733 32318 12767
rect 32505 12733 32539 12767
rect 32597 12665 32631 12699
rect 32413 12597 32447 12631
rect 2145 12393 2179 12427
rect 2053 12189 2087 12223
rect 67649 7837 67683 7871
rect 1869 7769 1903 7803
rect 67925 7769 67959 7803
rect 2145 7701 2179 7735
rect 67925 6749 67959 6783
rect 65809 6273 65843 6307
rect 65993 6205 66027 6239
rect 67557 6205 67591 6239
rect 67649 5865 67683 5899
rect 66453 5661 66487 5695
rect 66913 5661 66947 5695
rect 67557 5661 67591 5695
rect 67005 5525 67039 5559
rect 65993 5253 66027 5287
rect 65809 5117 65843 5151
rect 67557 5117 67591 5151
rect 6377 4641 6411 4675
rect 5641 4573 5675 4607
rect 66913 4573 66947 4607
rect 67373 4573 67407 4607
rect 67465 4437 67499 4471
rect 5089 4097 5123 4131
rect 6837 4097 6871 4131
rect 45753 4097 45787 4131
rect 61945 4097 61979 4131
rect 65809 4029 65843 4063
rect 65993 4029 66027 4063
rect 67649 4029 67683 4063
rect 1869 3893 1903 3927
rect 4629 3893 4663 3927
rect 5181 3893 5215 3927
rect 6929 3893 6963 3927
rect 45845 3893 45879 3927
rect 60933 3893 60967 3927
rect 62037 3893 62071 3927
rect 4445 3553 4479 3587
rect 4905 3553 4939 3587
rect 10977 3553 11011 3587
rect 46397 3553 46431 3587
rect 47041 3553 47075 3587
rect 62129 3553 62163 3587
rect 62497 3553 62531 3587
rect 1961 3485 1995 3519
rect 2789 3485 2823 3519
rect 6745 3485 6779 3519
rect 7573 3485 7607 3519
rect 10425 3485 10459 3519
rect 19625 3485 19659 3519
rect 22017 3485 22051 3519
rect 38393 3485 38427 3519
rect 45017 3485 45051 3519
rect 46213 3485 46247 3519
rect 60749 3485 60783 3519
rect 61945 3485 61979 3519
rect 67005 3485 67039 3519
rect 67465 3485 67499 3519
rect 4629 3417 4663 3451
rect 10609 3417 10643 3451
rect 2053 3349 2087 3383
rect 6837 3349 6871 3383
rect 22109 3349 22143 3383
rect 45109 3349 45143 3383
rect 60841 3349 60875 3383
rect 67557 3349 67591 3383
rect 1777 3077 1811 3111
rect 6837 3077 6871 3111
rect 10609 3077 10643 3111
rect 22109 3077 22143 3111
rect 33517 3077 33551 3111
rect 34253 3077 34287 3111
rect 44833 3077 44867 3111
rect 60841 3077 60875 3111
rect 65993 3077 66027 3111
rect 1593 3009 1627 3043
rect 3893 3009 3927 3043
rect 6653 3009 6687 3043
rect 10241 3009 10275 3043
rect 10517 3009 10551 3043
rect 19349 3009 19383 3043
rect 33425 3009 33459 3043
rect 38117 3009 38151 3043
rect 60657 3009 60691 3043
rect 65809 3009 65843 3043
rect 2789 2941 2823 2975
rect 4077 2941 4111 2975
rect 4353 2941 4387 2975
rect 7113 2941 7147 2975
rect 19533 2941 19567 2975
rect 19993 2941 20027 2975
rect 21925 2941 21959 2975
rect 22845 2941 22879 2975
rect 34069 2941 34103 2975
rect 34805 2941 34839 2975
rect 38301 2941 38335 2975
rect 38669 2941 38703 2975
rect 44189 2941 44223 2975
rect 44649 2941 44683 2975
rect 45109 2941 45143 2975
rect 61209 2941 61243 2975
rect 67649 2941 67683 2975
rect 2513 2601 2547 2635
rect 3985 2601 4019 2635
rect 10701 2601 10735 2635
rect 17693 2601 17727 2635
rect 19533 2601 19567 2635
rect 22753 2601 22787 2635
rect 32321 2601 32355 2635
rect 34897 2601 34931 2635
rect 38209 2601 38243 2635
rect 46397 2601 46431 2635
rect 62129 2601 62163 2635
rect 22017 2533 22051 2567
rect 43085 2533 43119 2567
rect 6561 2465 6595 2499
rect 6929 2465 6963 2499
rect 27445 2465 27479 2499
rect 2421 2397 2455 2431
rect 3801 2397 3835 2431
rect 5733 2397 5767 2431
rect 6377 2397 6411 2431
rect 17509 2397 17543 2431
rect 19441 2397 19475 2431
rect 21833 2397 21867 2431
rect 27169 2397 27203 2431
rect 28457 2397 28491 2431
rect 32505 2397 32539 2431
rect 38117 2397 38151 2431
rect 56149 2397 56183 2431
rect 65625 2397 65659 2431
rect 42901 2329 42935 2363
rect 56425 2329 56459 2363
rect 65901 2329 65935 2363
rect 67281 2329 67315 2363
rect 28641 2261 28675 2295
rect 67373 2261 67407 2295
<< metal1 >>
rect 1104 69658 68816 69680
rect 1104 69606 19574 69658
rect 19626 69606 19638 69658
rect 19690 69606 19702 69658
rect 19754 69606 19766 69658
rect 19818 69606 19830 69658
rect 19882 69606 50294 69658
rect 50346 69606 50358 69658
rect 50410 69606 50422 69658
rect 50474 69606 50486 69658
rect 50538 69606 50550 69658
rect 50602 69606 68816 69658
rect 1104 69584 68816 69606
rect 14182 69436 14188 69488
rect 14240 69476 14246 69488
rect 14553 69479 14611 69485
rect 14553 69476 14565 69479
rect 14240 69448 14565 69476
rect 14240 69436 14246 69448
rect 14553 69445 14565 69448
rect 14599 69445 14611 69479
rect 14553 69439 14611 69445
rect 19334 69436 19340 69488
rect 19392 69476 19398 69488
rect 19705 69479 19763 69485
rect 19705 69476 19717 69479
rect 19392 69448 19717 69476
rect 19392 69436 19398 69448
rect 19705 69445 19717 69448
rect 19751 69445 19763 69479
rect 19705 69439 19763 69445
rect 20622 69436 20628 69488
rect 20680 69476 20686 69488
rect 20809 69479 20867 69485
rect 20809 69476 20821 69479
rect 20680 69448 20821 69476
rect 20680 69436 20686 69448
rect 20809 69445 20821 69448
rect 20855 69445 20867 69479
rect 35618 69476 35624 69488
rect 35579 69448 35624 69476
rect 20809 69439 20867 69445
rect 35618 69436 35624 69448
rect 35676 69436 35682 69488
rect 67637 69479 67695 69485
rect 67637 69445 67649 69479
rect 67683 69476 67695 69479
rect 68278 69476 68284 69488
rect 67683 69448 68284 69476
rect 67683 69445 67695 69448
rect 67637 69439 67695 69445
rect 68278 69436 68284 69448
rect 68336 69436 68342 69488
rect 1394 69408 1400 69420
rect 1355 69380 1400 69408
rect 1394 69368 1400 69380
rect 1452 69368 1458 69420
rect 7742 69368 7748 69420
rect 7800 69408 7806 69420
rect 7837 69411 7895 69417
rect 7837 69408 7849 69411
rect 7800 69380 7849 69408
rect 7800 69368 7806 69380
rect 7837 69377 7849 69380
rect 7883 69377 7895 69411
rect 7837 69371 7895 69377
rect 46474 69368 46480 69420
rect 46532 69408 46538 69420
rect 46569 69411 46627 69417
rect 46569 69408 46581 69411
rect 46532 69380 46581 69408
rect 46532 69368 46538 69380
rect 46569 69377 46581 69380
rect 46615 69408 46627 69411
rect 46615 69380 55214 69408
rect 46615 69377 46627 69380
rect 46569 69371 46627 69377
rect 1578 69340 1584 69352
rect 1539 69312 1584 69340
rect 1578 69300 1584 69312
rect 1636 69300 1642 69352
rect 55186 69340 55214 69380
rect 55398 69368 55404 69420
rect 55456 69408 55462 69420
rect 55493 69411 55551 69417
rect 55493 69408 55505 69411
rect 55456 69380 55505 69408
rect 55456 69368 55462 69380
rect 55493 69377 55505 69380
rect 55539 69377 55551 69411
rect 55493 69371 55551 69377
rect 57238 69368 57244 69420
rect 57296 69408 57302 69420
rect 57885 69411 57943 69417
rect 57885 69408 57897 69411
rect 57296 69380 57897 69408
rect 57296 69368 57302 69380
rect 57885 69377 57897 69380
rect 57931 69377 57943 69411
rect 57885 69371 57943 69377
rect 59722 69340 59728 69352
rect 55186 69312 59728 69340
rect 59722 69300 59728 69312
rect 59780 69300 59786 69352
rect 65058 69300 65064 69352
rect 65116 69340 65122 69352
rect 65797 69343 65855 69349
rect 65797 69340 65809 69343
rect 65116 69312 65809 69340
rect 65116 69300 65122 69312
rect 65797 69309 65809 69312
rect 65843 69309 65855 69343
rect 65797 69303 65855 69309
rect 65981 69343 66039 69349
rect 65981 69309 65993 69343
rect 66027 69340 66039 69343
rect 66346 69340 66352 69352
rect 66027 69312 66352 69340
rect 66027 69309 66039 69312
rect 65981 69303 66039 69309
rect 66346 69300 66352 69312
rect 66404 69300 66410 69352
rect 14737 69275 14795 69281
rect 14737 69241 14749 69275
rect 14783 69272 14795 69275
rect 14826 69272 14832 69284
rect 14783 69244 14832 69272
rect 14783 69241 14795 69244
rect 14737 69235 14795 69241
rect 14826 69232 14832 69244
rect 14884 69232 14890 69284
rect 19889 69275 19947 69281
rect 19889 69241 19901 69275
rect 19935 69272 19947 69275
rect 20254 69272 20260 69284
rect 19935 69244 20260 69272
rect 19935 69241 19947 69244
rect 19889 69235 19947 69241
rect 20254 69232 20260 69244
rect 20312 69232 20318 69284
rect 20993 69275 21051 69281
rect 20993 69241 21005 69275
rect 21039 69272 21051 69275
rect 21634 69272 21640 69284
rect 21039 69244 21640 69272
rect 21039 69241 21051 69244
rect 20993 69235 21051 69241
rect 21634 69232 21640 69244
rect 21692 69232 21698 69284
rect 35897 69275 35955 69281
rect 35897 69241 35909 69275
rect 35943 69272 35955 69275
rect 36906 69272 36912 69284
rect 35943 69244 36912 69272
rect 35943 69241 35955 69244
rect 35897 69235 35955 69241
rect 36906 69232 36912 69244
rect 36964 69232 36970 69284
rect 2498 69204 2504 69216
rect 2459 69176 2504 69204
rect 2498 69164 2504 69176
rect 2556 69164 2562 69216
rect 4798 69204 4804 69216
rect 4759 69176 4804 69204
rect 4798 69164 4804 69176
rect 4856 69164 4862 69216
rect 5994 69164 6000 69216
rect 6052 69204 6058 69216
rect 6549 69207 6607 69213
rect 6549 69204 6561 69207
rect 6052 69176 6561 69204
rect 6052 69164 6058 69176
rect 6549 69173 6561 69176
rect 6595 69173 6607 69207
rect 8018 69204 8024 69216
rect 7979 69176 8024 69204
rect 6549 69167 6607 69173
rect 8018 69164 8024 69176
rect 8076 69164 8082 69216
rect 11698 69204 11704 69216
rect 11659 69176 11704 69204
rect 11698 69164 11704 69176
rect 11756 69164 11762 69216
rect 16850 69204 16856 69216
rect 16811 69176 16856 69204
rect 16850 69164 16856 69176
rect 16908 69164 16914 69216
rect 24854 69204 24860 69216
rect 24815 69176 24860 69204
rect 24854 69164 24860 69176
rect 24912 69164 24918 69216
rect 27338 69204 27344 69216
rect 27299 69176 27344 69204
rect 27338 69164 27344 69176
rect 27396 69164 27402 69216
rect 31202 69204 31208 69216
rect 31163 69176 31208 69204
rect 31202 69164 31208 69176
rect 31260 69164 31266 69216
rect 36630 69204 36636 69216
rect 36591 69176 36636 69204
rect 36630 69164 36636 69176
rect 36688 69164 36694 69216
rect 37274 69164 37280 69216
rect 37332 69204 37338 69216
rect 37553 69207 37611 69213
rect 37553 69204 37565 69207
rect 37332 69176 37565 69204
rect 37332 69164 37338 69176
rect 37553 69173 37565 69176
rect 37599 69173 37611 69207
rect 39022 69204 39028 69216
rect 38983 69176 39028 69204
rect 37553 69167 37611 69173
rect 39022 69164 39028 69176
rect 39080 69164 39086 69216
rect 41414 69204 41420 69216
rect 41375 69176 41420 69204
rect 41414 69164 41420 69176
rect 41472 69164 41478 69216
rect 42886 69204 42892 69216
rect 42847 69176 42892 69204
rect 42886 69164 42892 69176
rect 42944 69164 42950 69216
rect 45186 69164 45192 69216
rect 45244 69204 45250 69216
rect 45465 69207 45523 69213
rect 45465 69204 45477 69207
rect 45244 69176 45477 69204
rect 45244 69164 45250 69176
rect 45465 69173 45477 69176
rect 45511 69173 45523 69207
rect 46106 69204 46112 69216
rect 46067 69176 46112 69204
rect 45465 69167 45523 69173
rect 46106 69164 46112 69176
rect 46164 69164 46170 69216
rect 46566 69164 46572 69216
rect 46624 69204 46630 69216
rect 46661 69207 46719 69213
rect 46661 69204 46673 69207
rect 46624 69176 46673 69204
rect 46624 69164 46630 69176
rect 46661 69173 46673 69176
rect 46707 69173 46719 69207
rect 50706 69204 50712 69216
rect 50667 69176 50712 69204
rect 46661 69167 46719 69173
rect 50706 69164 50712 69176
rect 50764 69164 50770 69216
rect 52914 69204 52920 69216
rect 52875 69176 52920 69204
rect 52914 69164 52920 69176
rect 52972 69164 52978 69216
rect 55674 69204 55680 69216
rect 55635 69176 55680 69204
rect 55674 69164 55680 69176
rect 55732 69164 55738 69216
rect 56502 69204 56508 69216
rect 56463 69176 56508 69204
rect 56502 69164 56508 69176
rect 56560 69164 56566 69216
rect 57330 69204 57336 69216
rect 57291 69176 57336 69204
rect 57330 69164 57336 69176
rect 57388 69164 57394 69216
rect 57977 69207 58035 69213
rect 57977 69173 57989 69207
rect 58023 69204 58035 69207
rect 58066 69204 58072 69216
rect 58023 69176 58072 69204
rect 58023 69173 58035 69176
rect 57977 69167 58035 69173
rect 58066 69164 58072 69176
rect 58124 69164 58130 69216
rect 60642 69204 60648 69216
rect 60603 69176 60648 69204
rect 60642 69164 60648 69176
rect 60700 69164 60706 69216
rect 62206 69204 62212 69216
rect 62167 69176 62212 69204
rect 62206 69164 62212 69176
rect 62264 69164 62270 69216
rect 64417 69207 64475 69213
rect 64417 69173 64429 69207
rect 64463 69204 64475 69207
rect 64966 69204 64972 69216
rect 64463 69176 64972 69204
rect 64463 69173 64475 69176
rect 64417 69167 64475 69173
rect 64966 69164 64972 69176
rect 65024 69164 65030 69216
rect 65061 69207 65119 69213
rect 65061 69173 65073 69207
rect 65107 69204 65119 69207
rect 66254 69204 66260 69216
rect 65107 69176 66260 69204
rect 65107 69173 65119 69176
rect 65061 69167 65119 69173
rect 66254 69164 66260 69176
rect 66312 69164 66318 69216
rect 1104 69114 68816 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 34934 69114
rect 34986 69062 34998 69114
rect 35050 69062 35062 69114
rect 35114 69062 35126 69114
rect 35178 69062 35190 69114
rect 35242 69062 65654 69114
rect 65706 69062 65718 69114
rect 65770 69062 65782 69114
rect 65834 69062 65846 69114
rect 65898 69062 65910 69114
rect 65962 69062 68816 69114
rect 1104 69040 68816 69062
rect 11606 68892 11612 68944
rect 11664 68932 11670 68944
rect 11664 68904 11836 68932
rect 11664 68892 11670 68904
rect 1397 68867 1455 68873
rect 1397 68833 1409 68867
rect 1443 68864 1455 68867
rect 2498 68864 2504 68876
rect 1443 68836 2504 68864
rect 1443 68833 1455 68836
rect 1397 68827 1455 68833
rect 2498 68824 2504 68836
rect 2556 68824 2562 68876
rect 2774 68864 2780 68876
rect 2735 68836 2780 68864
rect 2774 68824 2780 68836
rect 2832 68824 2838 68876
rect 5994 68864 6000 68876
rect 5955 68836 6000 68864
rect 5994 68824 6000 68836
rect 6052 68824 6058 68876
rect 6454 68864 6460 68876
rect 6415 68836 6460 68864
rect 6454 68824 6460 68836
rect 6512 68824 6518 68876
rect 11057 68867 11115 68873
rect 11057 68833 11069 68867
rect 11103 68864 11115 68867
rect 11698 68864 11704 68876
rect 11103 68836 11704 68864
rect 11103 68833 11115 68836
rect 11057 68827 11115 68833
rect 11698 68824 11704 68836
rect 11756 68824 11762 68876
rect 11808 68873 11836 68904
rect 16758 68892 16764 68944
rect 16816 68932 16822 68944
rect 16816 68904 16988 68932
rect 16816 68892 16822 68904
rect 11793 68867 11851 68873
rect 11793 68833 11805 68867
rect 11839 68833 11851 68867
rect 11793 68827 11851 68833
rect 16117 68867 16175 68873
rect 16117 68833 16129 68867
rect 16163 68864 16175 68867
rect 16850 68864 16856 68876
rect 16163 68836 16856 68864
rect 16163 68833 16175 68836
rect 16117 68827 16175 68833
rect 16850 68824 16856 68836
rect 16908 68824 16914 68876
rect 16960 68873 16988 68904
rect 52822 68892 52828 68944
rect 52880 68932 52886 68944
rect 52880 68904 53236 68932
rect 52880 68892 52886 68904
rect 16945 68867 17003 68873
rect 16945 68833 16957 68867
rect 16991 68833 17003 68867
rect 16945 68827 17003 68833
rect 24673 68867 24731 68873
rect 24673 68833 24685 68867
rect 24719 68864 24731 68867
rect 24854 68864 24860 68876
rect 24719 68836 24860 68864
rect 24719 68833 24731 68836
rect 24673 68827 24731 68833
rect 24854 68824 24860 68836
rect 24912 68824 24918 68876
rect 25130 68864 25136 68876
rect 25091 68836 25136 68864
rect 25130 68824 25136 68836
rect 25188 68824 25194 68876
rect 27065 68867 27123 68873
rect 27065 68833 27077 68867
rect 27111 68864 27123 68867
rect 27338 68864 27344 68876
rect 27111 68836 27344 68864
rect 27111 68833 27123 68836
rect 27065 68827 27123 68833
rect 27338 68824 27344 68836
rect 27396 68824 27402 68876
rect 27706 68864 27712 68876
rect 27667 68836 27712 68864
rect 27706 68824 27712 68836
rect 27764 68824 27770 68876
rect 31021 68867 31079 68873
rect 31021 68833 31033 68867
rect 31067 68864 31079 68867
rect 31202 68864 31208 68876
rect 31067 68836 31208 68864
rect 31067 68833 31079 68836
rect 31021 68827 31079 68833
rect 31202 68824 31208 68836
rect 31260 68824 31266 68876
rect 31570 68824 31576 68876
rect 31628 68864 31634 68876
rect 31757 68867 31815 68873
rect 31757 68864 31769 68867
rect 31628 68836 31769 68864
rect 31628 68824 31634 68836
rect 31757 68833 31769 68836
rect 31803 68833 31815 68867
rect 31757 68827 31815 68833
rect 36265 68867 36323 68873
rect 36265 68833 36277 68867
rect 36311 68864 36323 68867
rect 36630 68864 36636 68876
rect 36311 68836 36636 68864
rect 36311 68833 36323 68836
rect 36265 68827 36323 68833
rect 36630 68824 36636 68836
rect 36688 68824 36694 68876
rect 36722 68824 36728 68876
rect 36780 68864 36786 68876
rect 40313 68867 40371 68873
rect 36780 68836 36825 68864
rect 36780 68824 36786 68836
rect 40313 68833 40325 68867
rect 40359 68864 40371 68867
rect 41414 68864 41420 68876
rect 40359 68836 41420 68864
rect 40359 68833 40371 68836
rect 40313 68827 40371 68833
rect 41414 68824 41420 68836
rect 41472 68824 41478 68876
rect 41874 68864 41880 68876
rect 41835 68836 41880 68864
rect 41874 68824 41880 68836
rect 41932 68824 41938 68876
rect 42613 68867 42671 68873
rect 42613 68833 42625 68867
rect 42659 68864 42671 68867
rect 42886 68864 42892 68876
rect 42659 68836 42892 68864
rect 42659 68833 42671 68836
rect 42613 68827 42671 68833
rect 42886 68824 42892 68836
rect 42944 68824 42950 68876
rect 43162 68864 43168 68876
rect 43123 68836 43168 68864
rect 43162 68824 43168 68836
rect 43220 68824 43226 68876
rect 46106 68824 46112 68876
rect 46164 68864 46170 68876
rect 46385 68867 46443 68873
rect 46385 68864 46397 68867
rect 46164 68836 46397 68864
rect 46164 68824 46170 68836
rect 46385 68833 46397 68836
rect 46431 68833 46443 68867
rect 46566 68864 46572 68876
rect 46527 68836 46572 68864
rect 46385 68827 46443 68833
rect 46566 68824 46572 68836
rect 46624 68824 46630 68876
rect 47026 68864 47032 68876
rect 46987 68836 47032 68864
rect 47026 68824 47032 68836
rect 47084 68824 47090 68876
rect 50433 68867 50491 68873
rect 50433 68833 50445 68867
rect 50479 68864 50491 68867
rect 50706 68864 50712 68876
rect 50479 68836 50712 68864
rect 50479 68833 50491 68836
rect 50433 68827 50491 68833
rect 50706 68824 50712 68836
rect 50764 68824 50770 68876
rect 51534 68864 51540 68876
rect 51495 68836 51540 68864
rect 51534 68824 51540 68836
rect 51592 68824 51598 68876
rect 52733 68867 52791 68873
rect 52733 68833 52745 68867
rect 52779 68864 52791 68867
rect 52914 68864 52920 68876
rect 52779 68836 52920 68864
rect 52779 68833 52791 68836
rect 52733 68827 52791 68833
rect 52914 68824 52920 68836
rect 52972 68824 52978 68876
rect 53208 68873 53236 68904
rect 60550 68892 60556 68944
rect 60608 68932 60614 68944
rect 60608 68904 60964 68932
rect 60608 68892 60614 68904
rect 53193 68867 53251 68873
rect 53193 68833 53205 68867
rect 53239 68833 53251 68867
rect 53193 68827 53251 68833
rect 56229 68867 56287 68873
rect 56229 68833 56241 68867
rect 56275 68864 56287 68867
rect 56502 68864 56508 68876
rect 56275 68836 56508 68864
rect 56275 68833 56287 68836
rect 56229 68827 56287 68833
rect 56502 68824 56508 68836
rect 56560 68824 56566 68876
rect 56686 68864 56692 68876
rect 56647 68836 56692 68864
rect 56686 68824 56692 68836
rect 56744 68824 56750 68876
rect 60461 68867 60519 68873
rect 60461 68833 60473 68867
rect 60507 68864 60519 68867
rect 60642 68864 60648 68876
rect 60507 68836 60648 68864
rect 60507 68833 60519 68836
rect 60461 68827 60519 68833
rect 60642 68824 60648 68836
rect 60700 68824 60706 68876
rect 60936 68873 60964 68904
rect 60921 68867 60979 68873
rect 60921 68833 60933 68867
rect 60967 68833 60979 68867
rect 60921 68827 60979 68833
rect 62206 68824 62212 68876
rect 62264 68864 62270 68876
rect 62761 68867 62819 68873
rect 62761 68864 62773 68867
rect 62264 68836 62773 68864
rect 62264 68824 62270 68836
rect 62761 68833 62773 68836
rect 62807 68833 62819 68867
rect 62761 68827 62819 68833
rect 63126 68824 63132 68876
rect 63184 68864 63190 68876
rect 63221 68867 63279 68873
rect 63221 68864 63233 68867
rect 63184 68836 63233 68864
rect 63184 68824 63190 68836
rect 63221 68833 63233 68836
rect 63267 68833 63279 68867
rect 66254 68864 66260 68876
rect 66215 68836 66260 68864
rect 63221 68827 63279 68833
rect 66254 68824 66260 68836
rect 66312 68824 66318 68876
rect 68097 68867 68155 68873
rect 68097 68833 68109 68867
rect 68143 68864 68155 68867
rect 69566 68864 69572 68876
rect 68143 68836 69572 68864
rect 68143 68833 68155 68836
rect 68097 68827 68155 68833
rect 69566 68824 69572 68836
rect 69624 68824 69630 68876
rect 4614 68796 4620 68808
rect 4575 68768 4620 68796
rect 4614 68756 4620 68768
rect 4672 68756 4678 68808
rect 5353 68799 5411 68805
rect 5353 68765 5365 68799
rect 5399 68796 5411 68799
rect 5902 68796 5908 68808
rect 5399 68768 5908 68796
rect 5399 68765 5411 68768
rect 5353 68759 5411 68765
rect 5902 68756 5908 68768
rect 5960 68756 5966 68808
rect 10410 68796 10416 68808
rect 10371 68768 10416 68796
rect 10410 68756 10416 68768
rect 10468 68756 10474 68808
rect 15470 68796 15476 68808
rect 15431 68768 15476 68796
rect 15470 68756 15476 68768
rect 15528 68756 15534 68808
rect 38930 68796 38936 68808
rect 38843 68768 38936 68796
rect 38930 68756 38936 68768
rect 38988 68796 38994 68808
rect 39850 68796 39856 68808
rect 38988 68768 39856 68796
rect 38988 68756 38994 68768
rect 39850 68756 39856 68768
rect 39908 68756 39914 68808
rect 45281 68799 45339 68805
rect 45281 68796 45293 68799
rect 44008 68768 45293 68796
rect 1581 68731 1639 68737
rect 1581 68697 1593 68731
rect 1627 68728 1639 68731
rect 1854 68728 1860 68740
rect 1627 68700 1860 68728
rect 1627 68697 1639 68700
rect 1581 68691 1639 68697
rect 1854 68688 1860 68700
rect 1912 68688 1918 68740
rect 5445 68731 5503 68737
rect 5445 68697 5457 68731
rect 5491 68728 5503 68731
rect 6181 68731 6239 68737
rect 6181 68728 6193 68731
rect 5491 68700 6193 68728
rect 5491 68697 5503 68700
rect 5445 68691 5503 68697
rect 6181 68697 6193 68700
rect 6227 68697 6239 68731
rect 6181 68691 6239 68697
rect 10505 68731 10563 68737
rect 10505 68697 10517 68731
rect 10551 68728 10563 68731
rect 11241 68731 11299 68737
rect 11241 68728 11253 68731
rect 10551 68700 11253 68728
rect 10551 68697 10563 68700
rect 10505 68691 10563 68697
rect 11241 68697 11253 68700
rect 11287 68697 11299 68731
rect 11241 68691 11299 68697
rect 15565 68731 15623 68737
rect 15565 68697 15577 68731
rect 15611 68728 15623 68731
rect 16301 68731 16359 68737
rect 16301 68728 16313 68731
rect 15611 68700 16313 68728
rect 15611 68697 15623 68700
rect 15565 68691 15623 68697
rect 16301 68697 16313 68700
rect 16347 68697 16359 68731
rect 24854 68728 24860 68740
rect 24815 68700 24860 68728
rect 16301 68691 16359 68697
rect 24854 68688 24860 68700
rect 24912 68688 24918 68740
rect 27246 68728 27252 68740
rect 27207 68700 27252 68728
rect 27246 68688 27252 68700
rect 27304 68688 27310 68740
rect 31202 68728 31208 68740
rect 31163 68700 31208 68728
rect 31202 68688 31208 68700
rect 31260 68688 31266 68740
rect 36449 68731 36507 68737
rect 36449 68697 36461 68731
rect 36495 68728 36507 68731
rect 36538 68728 36544 68740
rect 36495 68700 36544 68728
rect 36495 68697 36507 68700
rect 36449 68691 36507 68697
rect 36538 68688 36544 68700
rect 36596 68688 36602 68740
rect 40497 68731 40555 68737
rect 40497 68697 40509 68731
rect 40543 68728 40555 68731
rect 41414 68728 41420 68740
rect 40543 68700 41420 68728
rect 40543 68697 40555 68700
rect 40497 68691 40555 68697
rect 41414 68688 41420 68700
rect 41472 68688 41478 68740
rect 42794 68728 42800 68740
rect 42755 68700 42800 68728
rect 42794 68688 42800 68700
rect 42852 68688 42858 68740
rect 4706 68660 4712 68672
rect 4667 68632 4712 68660
rect 4706 68620 4712 68632
rect 4764 68620 4770 68672
rect 15470 68620 15476 68672
rect 15528 68660 15534 68672
rect 27154 68660 27160 68672
rect 15528 68632 27160 68660
rect 15528 68620 15534 68632
rect 27154 68620 27160 68632
rect 27212 68620 27218 68672
rect 39025 68663 39083 68669
rect 39025 68629 39037 68663
rect 39071 68660 39083 68663
rect 39758 68660 39764 68672
rect 39071 68632 39764 68660
rect 39071 68629 39083 68632
rect 39025 68623 39083 68629
rect 39758 68620 39764 68632
rect 39816 68620 39822 68672
rect 42610 68620 42616 68672
rect 42668 68660 42674 68672
rect 44008 68660 44036 68768
rect 45281 68765 45293 68768
rect 45327 68796 45339 68799
rect 48958 68796 48964 68808
rect 45327 68768 45554 68796
rect 48919 68768 48964 68796
rect 45327 68765 45339 68768
rect 45281 68759 45339 68765
rect 45526 68728 45554 68768
rect 48958 68756 48964 68768
rect 49016 68756 49022 68808
rect 49421 68799 49479 68805
rect 49421 68765 49433 68799
rect 49467 68765 49479 68799
rect 59722 68796 59728 68808
rect 59683 68768 59728 68796
rect 49421 68759 49479 68765
rect 49436 68728 49464 68759
rect 59722 68756 59728 68768
rect 59780 68756 59786 68808
rect 65613 68799 65671 68805
rect 65613 68796 65625 68799
rect 64846 68768 65625 68796
rect 45526 68700 49464 68728
rect 49513 68731 49571 68737
rect 49513 68697 49525 68731
rect 49559 68728 49571 68731
rect 50617 68731 50675 68737
rect 50617 68728 50629 68731
rect 49559 68700 50629 68728
rect 49559 68697 49571 68700
rect 49513 68691 49571 68697
rect 50617 68697 50629 68700
rect 50663 68697 50675 68731
rect 52914 68728 52920 68740
rect 52875 68700 52920 68728
rect 50617 68691 50675 68697
rect 52914 68688 52920 68700
rect 52972 68688 52978 68740
rect 56410 68728 56416 68740
rect 56371 68700 56416 68728
rect 56410 68688 56416 68700
rect 56468 68688 56474 68740
rect 59817 68731 59875 68737
rect 59817 68697 59829 68731
rect 59863 68728 59875 68731
rect 60645 68731 60703 68737
rect 60645 68728 60657 68731
rect 59863 68700 60657 68728
rect 59863 68697 59875 68700
rect 59817 68691 59875 68697
rect 60645 68697 60657 68700
rect 60691 68697 60703 68731
rect 62942 68728 62948 68740
rect 62903 68700 62948 68728
rect 60645 68691 60703 68697
rect 62942 68688 62948 68700
rect 63000 68688 63006 68740
rect 45370 68660 45376 68672
rect 42668 68632 44036 68660
rect 45331 68632 45376 68660
rect 42668 68620 42674 68632
rect 45370 68620 45376 68632
rect 45428 68620 45434 68672
rect 59722 68620 59728 68672
rect 59780 68660 59786 68672
rect 64846 68660 64874 68768
rect 65613 68765 65625 68768
rect 65659 68765 65671 68799
rect 65613 68759 65671 68765
rect 66441 68731 66499 68737
rect 66441 68697 66453 68731
rect 66487 68728 66499 68731
rect 67082 68728 67088 68740
rect 66487 68700 67088 68728
rect 66487 68697 66499 68700
rect 66441 68691 66499 68697
rect 67082 68688 67088 68700
rect 67140 68688 67146 68740
rect 65702 68660 65708 68672
rect 59780 68632 64874 68660
rect 65663 68632 65708 68660
rect 59780 68620 59786 68632
rect 65702 68620 65708 68632
rect 65760 68620 65766 68672
rect 1104 68570 68816 68592
rect 1104 68518 19574 68570
rect 19626 68518 19638 68570
rect 19690 68518 19702 68570
rect 19754 68518 19766 68570
rect 19818 68518 19830 68570
rect 19882 68518 50294 68570
rect 50346 68518 50358 68570
rect 50410 68518 50422 68570
rect 50474 68518 50486 68570
rect 50538 68518 50550 68570
rect 50602 68518 68816 68570
rect 1104 68496 68816 68518
rect 1854 68456 1860 68468
rect 1815 68428 1860 68456
rect 1854 68416 1860 68428
rect 1912 68416 1918 68468
rect 4614 68416 4620 68468
rect 4672 68456 4678 68468
rect 23290 68456 23296 68468
rect 4672 68428 23296 68456
rect 4672 68416 4678 68428
rect 23290 68416 23296 68428
rect 23348 68416 23354 68468
rect 24765 68459 24823 68465
rect 24765 68425 24777 68459
rect 24811 68456 24823 68459
rect 24854 68456 24860 68468
rect 24811 68428 24860 68456
rect 24811 68425 24823 68428
rect 24765 68419 24823 68425
rect 24854 68416 24860 68428
rect 24912 68416 24918 68468
rect 27246 68456 27252 68468
rect 27207 68428 27252 68456
rect 27246 68416 27252 68428
rect 27304 68416 27310 68468
rect 31113 68459 31171 68465
rect 31113 68425 31125 68459
rect 31159 68456 31171 68459
rect 31202 68456 31208 68468
rect 31159 68428 31208 68456
rect 31159 68425 31171 68428
rect 31113 68419 31171 68425
rect 31202 68416 31208 68428
rect 31260 68416 31266 68468
rect 36538 68456 36544 68468
rect 36499 68428 36544 68456
rect 36538 68416 36544 68428
rect 36596 68416 36602 68468
rect 42610 68456 42616 68468
rect 39592 68428 42616 68456
rect 39592 68388 39620 68428
rect 42610 68416 42616 68428
rect 42668 68416 42674 68468
rect 42794 68456 42800 68468
rect 42755 68428 42800 68456
rect 42794 68416 42800 68428
rect 42852 68416 42858 68468
rect 52825 68459 52883 68465
rect 42904 68428 45554 68456
rect 39758 68388 39764 68400
rect 29748 68360 39620 68388
rect 39719 68360 39764 68388
rect 1765 68323 1823 68329
rect 1765 68289 1777 68323
rect 1811 68289 1823 68323
rect 1765 68283 1823 68289
rect 1780 68252 1808 68283
rect 2038 68280 2044 68332
rect 2096 68320 2102 68332
rect 2501 68323 2559 68329
rect 2501 68320 2513 68323
rect 2096 68292 2513 68320
rect 2096 68280 2102 68292
rect 2501 68289 2513 68292
rect 2547 68289 2559 68323
rect 24670 68320 24676 68332
rect 24631 68292 24676 68320
rect 2501 68283 2559 68289
rect 24670 68280 24676 68292
rect 24728 68280 24734 68332
rect 27154 68320 27160 68332
rect 27067 68292 27160 68320
rect 27154 68280 27160 68292
rect 27212 68320 27218 68332
rect 29748 68320 29776 68360
rect 39758 68348 39764 68360
rect 39816 68348 39822 68400
rect 39850 68348 39856 68400
rect 39908 68388 39914 68400
rect 42904 68388 42932 68428
rect 45370 68388 45376 68400
rect 39908 68360 42932 68388
rect 45331 68360 45376 68388
rect 39908 68348 39914 68360
rect 45370 68348 45376 68360
rect 45428 68348 45434 68400
rect 45526 68388 45554 68428
rect 52825 68425 52837 68459
rect 52871 68456 52883 68459
rect 52914 68456 52920 68468
rect 52871 68428 52920 68456
rect 52871 68425 52883 68428
rect 52825 68419 52883 68425
rect 52914 68416 52920 68428
rect 52972 68416 52978 68468
rect 56321 68459 56379 68465
rect 56321 68425 56333 68459
rect 56367 68456 56379 68459
rect 56410 68456 56416 68468
rect 56367 68428 56416 68456
rect 56367 68425 56379 68428
rect 56321 68419 56379 68425
rect 56410 68416 56416 68428
rect 56468 68416 56474 68468
rect 61657 68459 61715 68465
rect 61657 68425 61669 68459
rect 61703 68456 61715 68459
rect 62942 68456 62948 68468
rect 61703 68428 62948 68456
rect 61703 68425 61715 68428
rect 61657 68419 61715 68425
rect 62942 68416 62948 68428
rect 63000 68416 63006 68468
rect 57238 68388 57244 68400
rect 45526 68360 57244 68388
rect 57238 68348 57244 68360
rect 57296 68348 57302 68400
rect 58066 68388 58072 68400
rect 58027 68360 58072 68388
rect 58066 68348 58072 68360
rect 58124 68348 58130 68400
rect 65702 68388 65708 68400
rect 65663 68360 65708 68388
rect 65702 68348 65708 68360
rect 65760 68348 65766 68400
rect 31018 68320 31024 68332
rect 27212 68292 29776 68320
rect 30979 68292 31024 68320
rect 27212 68280 27218 68292
rect 31018 68280 31024 68292
rect 31076 68280 31082 68332
rect 36446 68320 36452 68332
rect 36407 68292 36452 68320
rect 36446 68280 36452 68292
rect 36504 68280 36510 68332
rect 37274 68320 37280 68332
rect 37235 68292 37280 68320
rect 37274 68280 37280 68292
rect 37332 68280 37338 68332
rect 39022 68280 39028 68332
rect 39080 68320 39086 68332
rect 39577 68323 39635 68329
rect 39577 68320 39589 68323
rect 39080 68292 39589 68320
rect 39080 68280 39086 68292
rect 39577 68289 39589 68292
rect 39623 68289 39635 68323
rect 39577 68283 39635 68289
rect 42705 68323 42763 68329
rect 42705 68289 42717 68323
rect 42751 68289 42763 68323
rect 45186 68320 45192 68332
rect 45147 68292 45192 68320
rect 42705 68283 42763 68289
rect 3050 68252 3056 68264
rect 1780 68224 3056 68252
rect 3050 68212 3056 68224
rect 3108 68212 3114 68264
rect 3326 68252 3332 68264
rect 3287 68224 3332 68252
rect 3326 68212 3332 68224
rect 3384 68252 3390 68264
rect 37461 68255 37519 68261
rect 3384 68224 6914 68252
rect 3384 68212 3390 68224
rect 6886 68184 6914 68224
rect 37461 68221 37473 68255
rect 37507 68252 37519 68255
rect 37550 68252 37556 68264
rect 37507 68224 37556 68252
rect 37507 68221 37519 68224
rect 37461 68215 37519 68221
rect 37550 68212 37556 68224
rect 37608 68212 37614 68264
rect 38010 68252 38016 68264
rect 37971 68224 38016 68252
rect 38010 68212 38016 68224
rect 38068 68212 38074 68264
rect 39298 68212 39304 68264
rect 39356 68252 39362 68264
rect 40037 68255 40095 68261
rect 40037 68252 40049 68255
rect 39356 68224 40049 68252
rect 39356 68212 39362 68224
rect 40037 68221 40049 68224
rect 40083 68221 40095 68255
rect 40037 68215 40095 68221
rect 42720 68196 42748 68283
rect 45186 68280 45192 68292
rect 45244 68280 45250 68332
rect 48958 68280 48964 68332
rect 49016 68320 49022 68332
rect 49605 68323 49663 68329
rect 49605 68320 49617 68323
rect 49016 68292 49617 68320
rect 49016 68280 49022 68292
rect 49605 68289 49617 68292
rect 49651 68289 49663 68323
rect 52730 68320 52736 68332
rect 52691 68292 52736 68320
rect 49605 68283 49663 68289
rect 52730 68280 52736 68292
rect 52788 68280 52794 68332
rect 56226 68320 56232 68332
rect 56139 68292 56232 68320
rect 56226 68280 56232 68292
rect 56284 68320 56290 68332
rect 56284 68292 57284 68320
rect 56284 68280 56290 68292
rect 45738 68252 45744 68264
rect 45699 68224 45744 68252
rect 45738 68212 45744 68224
rect 45796 68212 45802 68264
rect 49789 68255 49847 68261
rect 49789 68221 49801 68255
rect 49835 68252 49847 68255
rect 50246 68252 50252 68264
rect 49835 68224 50252 68252
rect 49835 68221 49847 68224
rect 49789 68215 49847 68221
rect 50246 68212 50252 68224
rect 50304 68212 50310 68264
rect 50341 68255 50399 68261
rect 50341 68221 50353 68255
rect 50387 68221 50399 68255
rect 50341 68215 50399 68221
rect 42702 68184 42708 68196
rect 6886 68156 42708 68184
rect 42702 68144 42708 68156
rect 42760 68144 42766 68196
rect 50154 68144 50160 68196
rect 50212 68184 50218 68196
rect 50356 68184 50384 68215
rect 50212 68156 50384 68184
rect 57256 68184 57284 68292
rect 57330 68280 57336 68332
rect 57388 68320 57394 68332
rect 57885 68323 57943 68329
rect 57885 68320 57897 68323
rect 57388 68292 57897 68320
rect 57388 68280 57394 68292
rect 57885 68289 57897 68292
rect 57931 68289 57943 68323
rect 61562 68320 61568 68332
rect 61523 68292 61568 68320
rect 57885 68283 57943 68289
rect 61562 68280 61568 68292
rect 61620 68280 61626 68332
rect 64966 68280 64972 68332
rect 65024 68320 65030 68332
rect 65521 68323 65579 68329
rect 65521 68320 65533 68323
rect 65024 68292 65533 68320
rect 65024 68280 65030 68292
rect 65521 68289 65533 68292
rect 65567 68289 65579 68323
rect 65521 68283 65579 68289
rect 58066 68212 58072 68264
rect 58124 68252 58130 68264
rect 58345 68255 58403 68261
rect 58345 68252 58357 68255
rect 58124 68224 58357 68252
rect 58124 68212 58130 68224
rect 58345 68221 58357 68224
rect 58391 68221 58403 68255
rect 65058 68252 65064 68264
rect 65019 68224 65064 68252
rect 58345 68215 58403 68221
rect 65058 68212 65064 68224
rect 65116 68212 65122 68264
rect 66990 68252 66996 68264
rect 66951 68224 66996 68252
rect 66990 68212 66996 68224
rect 67048 68212 67054 68264
rect 67266 68184 67272 68196
rect 57256 68156 67272 68184
rect 50212 68144 50218 68156
rect 67266 68144 67272 68156
rect 67324 68144 67330 68196
rect 29178 68076 29184 68128
rect 29236 68116 29242 68128
rect 30282 68116 30288 68128
rect 29236 68088 30288 68116
rect 29236 68076 29242 68088
rect 30282 68076 30288 68088
rect 30340 68076 30346 68128
rect 1104 68026 68816 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 34934 68026
rect 34986 67974 34998 68026
rect 35050 67974 35062 68026
rect 35114 67974 35126 68026
rect 35178 67974 35190 68026
rect 35242 67974 65654 68026
rect 65706 67974 65718 68026
rect 65770 67974 65782 68026
rect 65834 67974 65846 68026
rect 65898 67974 65910 68026
rect 65962 67974 68816 68026
rect 1104 67952 68816 67974
rect 37550 67912 37556 67924
rect 37511 67884 37556 67912
rect 37550 67872 37556 67884
rect 37608 67872 37614 67924
rect 41414 67912 41420 67924
rect 41375 67884 41420 67912
rect 41414 67872 41420 67884
rect 41472 67872 41478 67924
rect 50246 67912 50252 67924
rect 50207 67884 50252 67912
rect 50246 67872 50252 67884
rect 50304 67872 50310 67924
rect 66257 67915 66315 67921
rect 66257 67881 66269 67915
rect 66303 67912 66315 67915
rect 66346 67912 66352 67924
rect 66303 67884 66352 67912
rect 66303 67881 66315 67884
rect 66257 67875 66315 67881
rect 66346 67872 66352 67884
rect 66404 67872 66410 67924
rect 67082 67912 67088 67924
rect 67043 67884 67088 67912
rect 67082 67872 67088 67884
rect 67140 67872 67146 67924
rect 4798 67844 4804 67856
rect 4540 67816 4804 67844
rect 2314 67776 2320 67788
rect 2275 67748 2320 67776
rect 2314 67736 2320 67748
rect 2372 67736 2378 67788
rect 4540 67785 4568 67816
rect 4798 67804 4804 67816
rect 4856 67804 4862 67856
rect 26206 67816 66760 67844
rect 4525 67779 4583 67785
rect 4525 67745 4537 67779
rect 4571 67745 4583 67779
rect 4706 67776 4712 67788
rect 4667 67748 4712 67776
rect 4525 67739 4583 67745
rect 4706 67736 4712 67748
rect 4764 67736 4770 67788
rect 5166 67776 5172 67788
rect 5127 67748 5172 67776
rect 5166 67736 5172 67748
rect 5224 67736 5230 67788
rect 24670 67776 24676 67788
rect 6886 67748 24676 67776
rect 2038 67708 2044 67720
rect 1999 67680 2044 67708
rect 2038 67668 2044 67680
rect 2096 67668 2102 67720
rect 2314 67600 2320 67652
rect 2372 67640 2378 67652
rect 6886 67640 6914 67748
rect 24670 67736 24676 67748
rect 24728 67776 24734 67788
rect 26206 67776 26234 67816
rect 24728 67748 26234 67776
rect 24728 67736 24734 67748
rect 31018 67736 31024 67788
rect 31076 67776 31082 67788
rect 31076 67748 55214 67776
rect 31076 67736 31082 67748
rect 37458 67708 37464 67720
rect 37419 67680 37464 67708
rect 37458 67668 37464 67680
rect 37516 67668 37522 67720
rect 41322 67708 41328 67720
rect 41283 67680 41328 67708
rect 41322 67668 41328 67680
rect 41380 67668 41386 67720
rect 50154 67708 50160 67720
rect 50115 67680 50160 67708
rect 50154 67668 50160 67680
rect 50212 67668 50218 67720
rect 55186 67708 55214 67748
rect 66732 67720 66760 67816
rect 66165 67711 66223 67717
rect 66165 67708 66177 67711
rect 55186 67680 66177 67708
rect 66165 67677 66177 67680
rect 66211 67677 66223 67711
rect 66165 67671 66223 67677
rect 66714 67668 66720 67720
rect 66772 67708 66778 67720
rect 66993 67711 67051 67717
rect 66993 67708 67005 67711
rect 66772 67680 67005 67708
rect 66772 67668 66778 67680
rect 66993 67677 67005 67680
rect 67039 67677 67051 67711
rect 67726 67708 67732 67720
rect 67687 67680 67732 67708
rect 66993 67671 67051 67677
rect 67726 67668 67732 67680
rect 67784 67668 67790 67720
rect 2372 67612 6914 67640
rect 2372 67600 2378 67612
rect 38562 67600 38568 67652
rect 38620 67640 38626 67652
rect 68097 67643 68155 67649
rect 68097 67640 68109 67643
rect 38620 67612 68109 67640
rect 38620 67600 38626 67612
rect 68097 67609 68109 67612
rect 68143 67609 68155 67643
rect 68097 67603 68155 67609
rect 1104 67482 68816 67504
rect 1104 67430 19574 67482
rect 19626 67430 19638 67482
rect 19690 67430 19702 67482
rect 19754 67430 19766 67482
rect 19818 67430 19830 67482
rect 19882 67430 50294 67482
rect 50346 67430 50358 67482
rect 50410 67430 50422 67482
rect 50474 67430 50486 67482
rect 50538 67430 50550 67482
rect 50602 67430 68816 67482
rect 1104 67408 68816 67430
rect 67634 67300 67640 67312
rect 67595 67272 67640 67300
rect 67634 67260 67640 67272
rect 67692 67260 67698 67312
rect 1578 67232 1584 67244
rect 1491 67204 1584 67232
rect 1578 67192 1584 67204
rect 1636 67192 1642 67244
rect 1857 67235 1915 67241
rect 1857 67201 1869 67235
rect 1903 67232 1915 67235
rect 2038 67232 2044 67244
rect 1903 67204 2044 67232
rect 1903 67201 1915 67204
rect 1857 67195 1915 67201
rect 2038 67192 2044 67204
rect 2096 67232 2102 67244
rect 2590 67232 2596 67244
rect 2096 67204 2596 67232
rect 2096 67192 2102 67204
rect 2590 67192 2596 67204
rect 2648 67232 2654 67244
rect 2685 67235 2743 67241
rect 2685 67232 2697 67235
rect 2648 67204 2697 67232
rect 2648 67192 2654 67204
rect 2685 67201 2697 67204
rect 2731 67232 2743 67235
rect 4341 67235 4399 67241
rect 4341 67232 4353 67235
rect 2731 67204 4353 67232
rect 2731 67201 2743 67204
rect 2685 67195 2743 67201
rect 4341 67201 4353 67204
rect 4387 67201 4399 67235
rect 4341 67195 4399 67201
rect 1596 67164 1624 67192
rect 2866 67164 2872 67176
rect 1596 67136 2872 67164
rect 2866 67124 2872 67136
rect 2924 67124 2930 67176
rect 3050 67164 3056 67176
rect 3011 67136 3056 67164
rect 3050 67124 3056 67136
rect 3108 67124 3114 67176
rect 5166 67164 5172 67176
rect 5127 67136 5172 67164
rect 5166 67124 5172 67136
rect 5224 67164 5230 67176
rect 40954 67164 40960 67176
rect 5224 67136 40960 67164
rect 5224 67124 5230 67136
rect 40954 67124 40960 67136
rect 41012 67164 41018 67176
rect 41322 67164 41328 67176
rect 41012 67136 41328 67164
rect 41012 67124 41018 67136
rect 41322 67124 41328 67136
rect 41380 67124 41386 67176
rect 65797 67167 65855 67173
rect 65797 67133 65809 67167
rect 65843 67133 65855 67167
rect 65797 67127 65855 67133
rect 65981 67167 66039 67173
rect 65981 67133 65993 67167
rect 66027 67164 66039 67167
rect 67542 67164 67548 67176
rect 66027 67136 67548 67164
rect 66027 67133 66039 67136
rect 65981 67127 66039 67133
rect 3068 67096 3096 67124
rect 36446 67096 36452 67108
rect 3068 67068 36452 67096
rect 36446 67056 36452 67068
rect 36504 67096 36510 67108
rect 36998 67096 37004 67108
rect 36504 67068 37004 67096
rect 36504 67056 36510 67068
rect 36998 67056 37004 67068
rect 37056 67056 37062 67108
rect 65812 67096 65840 67127
rect 67542 67124 67548 67136
rect 67600 67124 67606 67176
rect 66990 67096 66996 67108
rect 65812 67068 66996 67096
rect 66990 67056 66996 67068
rect 67048 67056 67054 67108
rect 1104 66938 68816 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 34934 66938
rect 34986 66886 34998 66938
rect 35050 66886 35062 66938
rect 35114 66886 35126 66938
rect 35178 66886 35190 66938
rect 35242 66886 65654 66938
rect 65706 66886 65718 66938
rect 65770 66886 65782 66938
rect 65834 66886 65846 66938
rect 65898 66886 65910 66938
rect 65962 66886 68816 66938
rect 1104 66864 68816 66886
rect 66990 66824 66996 66836
rect 66951 66796 66996 66824
rect 66990 66784 66996 66796
rect 67048 66784 67054 66836
rect 67542 66824 67548 66836
rect 67503 66796 67548 66824
rect 67542 66784 67548 66796
rect 67600 66784 67606 66836
rect 2774 66688 2780 66700
rect 2735 66660 2780 66688
rect 2774 66648 2780 66660
rect 2832 66648 2838 66700
rect 5902 66648 5908 66700
rect 5960 66688 5966 66700
rect 5997 66691 6055 66697
rect 5997 66688 6009 66691
rect 5960 66660 6009 66688
rect 5960 66648 5966 66660
rect 5997 66657 6009 66660
rect 6043 66688 6055 66691
rect 10410 66688 10416 66700
rect 6043 66660 10416 66688
rect 6043 66657 6055 66660
rect 5997 66651 6055 66657
rect 10410 66648 10416 66660
rect 10468 66648 10474 66700
rect 1394 66620 1400 66632
rect 1355 66592 1400 66620
rect 1394 66580 1400 66592
rect 1452 66580 1458 66632
rect 3973 66623 4031 66629
rect 3973 66589 3985 66623
rect 4019 66620 4031 66623
rect 4062 66620 4068 66632
rect 4019 66592 4068 66620
rect 4019 66589 4031 66592
rect 3973 66583 4031 66589
rect 4062 66580 4068 66592
rect 4120 66620 4126 66632
rect 5629 66623 5687 66629
rect 5629 66620 5641 66623
rect 4120 66592 5641 66620
rect 4120 66580 4126 66592
rect 5629 66589 5641 66592
rect 5675 66589 5687 66623
rect 5629 66583 5687 66589
rect 50154 66580 50160 66632
rect 50212 66620 50218 66632
rect 67450 66620 67456 66632
rect 50212 66592 67456 66620
rect 50212 66580 50218 66592
rect 67450 66580 67456 66592
rect 67508 66580 67514 66632
rect 1578 66552 1584 66564
rect 1539 66524 1584 66552
rect 1578 66512 1584 66524
rect 1636 66512 1642 66564
rect 4985 66555 5043 66561
rect 4985 66521 4997 66555
rect 5031 66521 5043 66555
rect 4985 66515 5043 66521
rect 4706 66444 4712 66496
rect 4764 66484 4770 66496
rect 5000 66484 5028 66515
rect 37458 66484 37464 66496
rect 4764 66456 37464 66484
rect 4764 66444 4770 66456
rect 37458 66444 37464 66456
rect 37516 66444 37522 66496
rect 1104 66394 68816 66416
rect 1104 66342 19574 66394
rect 19626 66342 19638 66394
rect 19690 66342 19702 66394
rect 19754 66342 19766 66394
rect 19818 66342 19830 66394
rect 19882 66342 50294 66394
rect 50346 66342 50358 66394
rect 50410 66342 50422 66394
rect 50474 66342 50486 66394
rect 50538 66342 50550 66394
rect 50602 66342 68816 66394
rect 1104 66320 68816 66342
rect 1578 66240 1584 66292
rect 1636 66280 1642 66292
rect 1949 66283 2007 66289
rect 1949 66280 1961 66283
rect 1636 66252 1961 66280
rect 1636 66240 1642 66252
rect 1949 66249 1961 66252
rect 1995 66249 2007 66283
rect 1949 66243 2007 66249
rect 1872 66184 6914 66212
rect 1872 66153 1900 66184
rect 1857 66147 1915 66153
rect 1857 66113 1869 66147
rect 1903 66113 1915 66147
rect 2590 66144 2596 66156
rect 2551 66116 2596 66144
rect 1857 66107 1915 66113
rect 2590 66104 2596 66116
rect 2648 66104 2654 66156
rect 4062 66104 4068 66156
rect 4120 66144 4126 66156
rect 4341 66147 4399 66153
rect 4341 66144 4353 66147
rect 4120 66116 4353 66144
rect 4120 66104 4126 66116
rect 4341 66113 4353 66116
rect 4387 66113 4399 66147
rect 6886 66144 6914 66184
rect 25130 66144 25136 66156
rect 6886 66116 25136 66144
rect 4341 66107 4399 66113
rect 25130 66104 25136 66116
rect 25188 66104 25194 66156
rect 36078 66144 36084 66156
rect 36039 66116 36084 66144
rect 36078 66104 36084 66116
rect 36136 66104 36142 66156
rect 52730 66144 52736 66156
rect 36280 66116 52736 66144
rect 3697 66079 3755 66085
rect 3697 66045 3709 66079
rect 3743 66045 3755 66079
rect 3697 66039 3755 66045
rect 3418 65968 3424 66020
rect 3476 66008 3482 66020
rect 3712 66008 3740 66039
rect 5258 66036 5264 66088
rect 5316 66076 5322 66088
rect 5537 66079 5595 66085
rect 5537 66076 5549 66079
rect 5316 66048 5549 66076
rect 5316 66036 5322 66048
rect 5537 66045 5549 66048
rect 5583 66076 5595 66079
rect 36280 66076 36308 66116
rect 52730 66104 52736 66116
rect 52788 66144 52794 66156
rect 53098 66144 53104 66156
rect 52788 66116 53104 66144
rect 52788 66104 52794 66116
rect 53098 66104 53104 66116
rect 53156 66104 53162 66156
rect 5583 66048 36308 66076
rect 5583 66045 5595 66048
rect 5537 66039 5595 66045
rect 36354 66036 36360 66088
rect 36412 66076 36418 66088
rect 65797 66079 65855 66085
rect 36412 66048 36457 66076
rect 36412 66036 36418 66048
rect 65797 66045 65809 66079
rect 65843 66045 65855 66079
rect 65797 66039 65855 66045
rect 65981 66079 66039 66085
rect 65981 66045 65993 66079
rect 66027 66076 66039 66079
rect 67358 66076 67364 66088
rect 66027 66048 67364 66076
rect 66027 66045 66039 66048
rect 65981 66039 66039 66045
rect 46474 66008 46480 66020
rect 3476 65980 46480 66008
rect 3476 65968 3482 65980
rect 46474 65968 46480 65980
rect 46532 65968 46538 66020
rect 65812 66008 65840 66039
rect 67358 66036 67364 66048
rect 67416 66036 67422 66088
rect 67542 66076 67548 66088
rect 67503 66048 67548 66076
rect 67542 66036 67548 66048
rect 67600 66036 67606 66088
rect 66990 66008 66996 66020
rect 65812 65980 66996 66008
rect 66990 65968 66996 65980
rect 67048 65968 67054 66020
rect 35894 65900 35900 65952
rect 35952 65940 35958 65952
rect 36265 65943 36323 65949
rect 35952 65912 35997 65940
rect 35952 65900 35958 65912
rect 36265 65909 36277 65943
rect 36311 65940 36323 65943
rect 36354 65940 36360 65952
rect 36311 65912 36360 65940
rect 36311 65909 36323 65912
rect 36265 65903 36323 65909
rect 36354 65900 36360 65912
rect 36412 65900 36418 65952
rect 1104 65850 68816 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 34934 65850
rect 34986 65798 34998 65850
rect 35050 65798 35062 65850
rect 35114 65798 35126 65850
rect 35178 65798 35190 65850
rect 35242 65798 65654 65850
rect 65706 65798 65718 65850
rect 65770 65798 65782 65850
rect 65834 65798 65846 65850
rect 65898 65798 65910 65850
rect 65962 65798 68816 65850
rect 1104 65776 68816 65798
rect 66990 65736 66996 65748
rect 66951 65708 66996 65736
rect 66990 65696 66996 65708
rect 67048 65696 67054 65748
rect 67358 65696 67364 65748
rect 67416 65736 67422 65748
rect 67545 65739 67603 65745
rect 67545 65736 67557 65739
rect 67416 65708 67557 65736
rect 67416 65696 67422 65708
rect 67545 65705 67557 65708
rect 67591 65705 67603 65739
rect 67545 65699 67603 65705
rect 1673 65535 1731 65541
rect 1673 65501 1685 65535
rect 1719 65532 1731 65535
rect 1762 65532 1768 65544
rect 1719 65504 1768 65532
rect 1719 65501 1731 65504
rect 1673 65495 1731 65501
rect 1762 65492 1768 65504
rect 1820 65492 1826 65544
rect 2133 65535 2191 65541
rect 2133 65501 2145 65535
rect 2179 65532 2191 65535
rect 3237 65535 3295 65541
rect 2179 65504 3188 65532
rect 2179 65501 2191 65504
rect 2133 65495 2191 65501
rect 2866 65464 2872 65476
rect 2779 65436 2872 65464
rect 2866 65424 2872 65436
rect 2924 65424 2930 65476
rect 3160 65464 3188 65504
rect 3237 65501 3249 65535
rect 3283 65532 3295 65535
rect 3973 65535 4031 65541
rect 3973 65532 3985 65535
rect 3283 65504 3985 65532
rect 3283 65501 3295 65504
rect 3237 65495 3295 65501
rect 3973 65501 3985 65504
rect 4019 65532 4031 65535
rect 4062 65532 4068 65544
rect 4019 65504 4068 65532
rect 4019 65501 4031 65504
rect 3973 65495 4031 65501
rect 4062 65492 4068 65504
rect 4120 65492 4126 65544
rect 33962 65492 33968 65544
rect 34020 65532 34026 65544
rect 35161 65535 35219 65541
rect 35161 65532 35173 65535
rect 34020 65504 35173 65532
rect 34020 65492 34026 65504
rect 35161 65501 35173 65504
rect 35207 65501 35219 65535
rect 35161 65495 35219 65501
rect 35428 65535 35486 65541
rect 35428 65501 35440 65535
rect 35474 65532 35486 65535
rect 35894 65532 35900 65544
rect 35474 65504 35900 65532
rect 35474 65501 35486 65504
rect 35428 65495 35486 65501
rect 35894 65492 35900 65504
rect 35952 65492 35958 65544
rect 67266 65492 67272 65544
rect 67324 65532 67330 65544
rect 67453 65535 67511 65541
rect 67453 65532 67465 65535
rect 67324 65504 67465 65532
rect 67324 65492 67330 65504
rect 67453 65501 67465 65504
rect 67499 65501 67511 65535
rect 67453 65495 67511 65501
rect 4338 65464 4344 65476
rect 3160 65436 4344 65464
rect 4338 65424 4344 65436
rect 4396 65424 4402 65476
rect 4798 65464 4804 65476
rect 4759 65436 4804 65464
rect 4798 65424 4804 65436
rect 4856 65424 4862 65476
rect 1946 65356 1952 65408
rect 2004 65396 2010 65408
rect 2225 65399 2283 65405
rect 2225 65396 2237 65399
rect 2004 65368 2237 65396
rect 2004 65356 2010 65368
rect 2225 65365 2237 65368
rect 2271 65365 2283 65399
rect 2884 65396 2912 65424
rect 23106 65396 23112 65408
rect 2884 65368 23112 65396
rect 2225 65359 2283 65365
rect 23106 65356 23112 65368
rect 23164 65356 23170 65408
rect 36262 65356 36268 65408
rect 36320 65396 36326 65408
rect 36541 65399 36599 65405
rect 36541 65396 36553 65399
rect 36320 65368 36553 65396
rect 36320 65356 36326 65368
rect 36541 65365 36553 65368
rect 36587 65365 36599 65399
rect 36541 65359 36599 65365
rect 1104 65306 68816 65328
rect 1104 65254 19574 65306
rect 19626 65254 19638 65306
rect 19690 65254 19702 65306
rect 19754 65254 19766 65306
rect 19818 65254 19830 65306
rect 19882 65254 50294 65306
rect 50346 65254 50358 65306
rect 50410 65254 50422 65306
rect 50474 65254 50486 65306
rect 50538 65254 50550 65306
rect 50602 65254 68816 65306
rect 1104 65232 68816 65254
rect 4798 65152 4804 65204
rect 4856 65192 4862 65204
rect 50154 65192 50160 65204
rect 4856 65164 50160 65192
rect 4856 65152 4862 65164
rect 50154 65152 50160 65164
rect 50212 65152 50218 65204
rect 1946 65124 1952 65136
rect 1907 65096 1952 65124
rect 1946 65084 1952 65096
rect 2004 65084 2010 65136
rect 1762 65056 1768 65068
rect 1723 65028 1768 65056
rect 1762 65016 1768 65028
rect 1820 65016 1826 65068
rect 4062 65056 4068 65068
rect 4023 65028 4068 65056
rect 4062 65016 4068 65028
rect 4120 65016 4126 65068
rect 36078 65056 36084 65068
rect 36039 65028 36084 65056
rect 36078 65016 36084 65028
rect 36136 65016 36142 65068
rect 36262 65056 36268 65068
rect 36223 65028 36268 65056
rect 36262 65016 36268 65028
rect 36320 65016 36326 65068
rect 36354 65016 36360 65068
rect 36412 65056 36418 65068
rect 38286 65056 38292 65068
rect 36412 65028 36457 65056
rect 38247 65028 38292 65056
rect 36412 65016 36418 65028
rect 38286 65016 38292 65028
rect 38344 65016 38350 65068
rect 3602 64988 3608 65000
rect 3563 64960 3608 64988
rect 3602 64948 3608 64960
rect 3660 64948 3666 65000
rect 4338 64988 4344 65000
rect 4251 64960 4344 64988
rect 4338 64948 4344 64960
rect 4396 64988 4402 65000
rect 15470 64988 15476 65000
rect 4396 64960 15476 64988
rect 4396 64948 4402 64960
rect 15470 64948 15476 64960
rect 15528 64948 15534 65000
rect 35897 64991 35955 64997
rect 35897 64957 35909 64991
rect 35943 64988 35955 64991
rect 36538 64988 36544 65000
rect 35943 64960 36544 64988
rect 35943 64957 35955 64960
rect 35897 64951 35955 64957
rect 36538 64948 36544 64960
rect 36596 64948 36602 65000
rect 38105 64855 38163 64861
rect 38105 64821 38117 64855
rect 38151 64852 38163 64855
rect 38194 64852 38200 64864
rect 38151 64824 38200 64852
rect 38151 64821 38163 64824
rect 38105 64815 38163 64821
rect 38194 64812 38200 64824
rect 38252 64812 38258 64864
rect 1104 64762 68816 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 34934 64762
rect 34986 64710 34998 64762
rect 35050 64710 35062 64762
rect 35114 64710 35126 64762
rect 35178 64710 35190 64762
rect 35242 64710 65654 64762
rect 65706 64710 65718 64762
rect 65770 64710 65782 64762
rect 65834 64710 65846 64762
rect 65898 64710 65910 64762
rect 65962 64710 68816 64762
rect 1104 64688 68816 64710
rect 1394 64608 1400 64660
rect 1452 64648 1458 64660
rect 1949 64651 2007 64657
rect 1949 64648 1961 64651
rect 1452 64620 1961 64648
rect 1452 64608 1458 64620
rect 1949 64617 1961 64620
rect 1995 64617 2007 64651
rect 1949 64611 2007 64617
rect 37277 64651 37335 64657
rect 37277 64617 37289 64651
rect 37323 64617 37335 64651
rect 37277 64611 37335 64617
rect 37461 64651 37519 64657
rect 37461 64617 37473 64651
rect 37507 64648 37519 64651
rect 38286 64648 38292 64660
rect 37507 64620 38292 64648
rect 37507 64617 37519 64620
rect 37461 64611 37519 64617
rect 36354 64540 36360 64592
rect 36412 64580 36418 64592
rect 36722 64580 36728 64592
rect 36412 64552 36728 64580
rect 36412 64540 36418 64552
rect 36722 64540 36728 64552
rect 36780 64580 36786 64592
rect 36909 64583 36967 64589
rect 36909 64580 36921 64583
rect 36780 64552 36921 64580
rect 36780 64540 36786 64552
rect 36909 64549 36921 64552
rect 36955 64549 36967 64583
rect 36909 64543 36967 64549
rect 36265 64447 36323 64453
rect 36265 64413 36277 64447
rect 36311 64444 36323 64447
rect 36630 64444 36636 64456
rect 36311 64416 36636 64444
rect 36311 64413 36323 64416
rect 36265 64407 36323 64413
rect 36630 64404 36636 64416
rect 36688 64444 36694 64456
rect 37292 64444 37320 64611
rect 38286 64608 38292 64620
rect 38344 64608 38350 64660
rect 38194 64453 38200 64456
rect 36688 64416 37320 64444
rect 37921 64447 37979 64453
rect 36688 64404 36694 64416
rect 37921 64413 37933 64447
rect 37967 64444 37979 64447
rect 37967 64416 38148 64444
rect 37967 64413 37979 64416
rect 37921 64407 37979 64413
rect 38120 64388 38148 64416
rect 38188 64407 38200 64453
rect 38252 64444 38258 64456
rect 38252 64416 38288 64444
rect 38194 64404 38200 64407
rect 38252 64404 38258 64416
rect 36449 64379 36507 64385
rect 36449 64345 36461 64379
rect 36495 64376 36507 64379
rect 36538 64376 36544 64388
rect 36495 64348 36544 64376
rect 36495 64345 36507 64348
rect 36449 64339 36507 64345
rect 36538 64336 36544 64348
rect 36596 64336 36602 64388
rect 38102 64336 38108 64388
rect 38160 64336 38166 64388
rect 37274 64308 37280 64320
rect 37235 64280 37280 64308
rect 37274 64268 37280 64280
rect 37332 64268 37338 64320
rect 37734 64268 37740 64320
rect 37792 64308 37798 64320
rect 39301 64311 39359 64317
rect 39301 64308 39313 64311
rect 37792 64280 39313 64308
rect 37792 64268 37798 64280
rect 39301 64277 39313 64280
rect 39347 64277 39359 64311
rect 39301 64271 39359 64277
rect 1104 64218 68816 64240
rect 1104 64166 19574 64218
rect 19626 64166 19638 64218
rect 19690 64166 19702 64218
rect 19754 64166 19766 64218
rect 19818 64166 19830 64218
rect 19882 64166 50294 64218
rect 50346 64166 50358 64218
rect 50410 64166 50422 64218
rect 50474 64166 50486 64218
rect 50538 64166 50550 64218
rect 50602 64166 68816 64218
rect 1104 64144 68816 64166
rect 36722 64104 36728 64116
rect 36683 64076 36728 64104
rect 36722 64064 36728 64076
rect 36780 64064 36786 64116
rect 37274 64064 37280 64116
rect 37332 64104 37338 64116
rect 37553 64107 37611 64113
rect 37553 64104 37565 64107
rect 37332 64076 37565 64104
rect 37332 64064 37338 64076
rect 37553 64073 37565 64076
rect 37599 64073 37611 64107
rect 37553 64067 37611 64073
rect 37921 64107 37979 64113
rect 37921 64073 37933 64107
rect 37967 64104 37979 64107
rect 38010 64104 38016 64116
rect 37967 64076 38016 64104
rect 37967 64073 37979 64076
rect 37921 64067 37979 64073
rect 38010 64064 38016 64076
rect 38068 64064 38074 64116
rect 36357 64039 36415 64045
rect 36357 64005 36369 64039
rect 36403 64005 36415 64039
rect 36357 63999 36415 64005
rect 36573 64039 36631 64045
rect 36573 64005 36585 64039
rect 36619 64036 36631 64039
rect 37642 64036 37648 64048
rect 36619 64008 37648 64036
rect 36619 64005 36631 64008
rect 36573 63999 36631 64005
rect 34232 63971 34290 63977
rect 34232 63937 34244 63971
rect 34278 63968 34290 63971
rect 34698 63968 34704 63980
rect 34278 63940 34704 63968
rect 34278 63937 34290 63940
rect 34232 63931 34290 63937
rect 34698 63928 34704 63940
rect 34756 63928 34762 63980
rect 36372 63968 36400 63999
rect 37642 63996 37648 64008
rect 37700 63996 37706 64048
rect 36814 63968 36820 63980
rect 36372 63940 36820 63968
rect 36814 63928 36820 63940
rect 36872 63968 36878 63980
rect 37734 63968 37740 63980
rect 36872 63940 37740 63968
rect 36872 63928 36878 63940
rect 37734 63928 37740 63940
rect 37792 63928 37798 63980
rect 38013 63971 38071 63977
rect 38013 63937 38025 63971
rect 38059 63937 38071 63971
rect 38013 63931 38071 63937
rect 33410 63860 33416 63912
rect 33468 63900 33474 63912
rect 33962 63900 33968 63912
rect 33468 63872 33968 63900
rect 33468 63860 33474 63872
rect 33962 63860 33968 63872
rect 34020 63860 34026 63912
rect 37642 63860 37648 63912
rect 37700 63900 37706 63912
rect 38028 63900 38056 63931
rect 37700 63872 38056 63900
rect 37700 63860 37706 63872
rect 35342 63764 35348 63776
rect 35303 63736 35348 63764
rect 35342 63724 35348 63736
rect 35400 63724 35406 63776
rect 36541 63767 36599 63773
rect 36541 63733 36553 63767
rect 36587 63764 36599 63767
rect 37274 63764 37280 63776
rect 36587 63736 37280 63764
rect 36587 63733 36599 63736
rect 36541 63727 36599 63733
rect 37274 63724 37280 63736
rect 37332 63724 37338 63776
rect 66254 63724 66260 63776
rect 66312 63764 66318 63776
rect 67637 63767 67695 63773
rect 67637 63764 67649 63767
rect 66312 63736 67649 63764
rect 66312 63724 66318 63736
rect 67637 63733 67649 63736
rect 67683 63733 67695 63767
rect 67637 63727 67695 63733
rect 1104 63674 68816 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 34934 63674
rect 34986 63622 34998 63674
rect 35050 63622 35062 63674
rect 35114 63622 35126 63674
rect 35178 63622 35190 63674
rect 35242 63622 65654 63674
rect 65706 63622 65718 63674
rect 65770 63622 65782 63674
rect 65834 63622 65846 63674
rect 65898 63622 65910 63674
rect 65962 63622 68816 63674
rect 1104 63600 68816 63622
rect 34698 63560 34704 63572
rect 34659 63532 34704 63560
rect 34698 63520 34704 63532
rect 34756 63520 34762 63572
rect 35802 63520 35808 63572
rect 35860 63560 35866 63572
rect 35989 63563 36047 63569
rect 35989 63560 36001 63563
rect 35860 63532 36001 63560
rect 35860 63520 35866 63532
rect 35989 63529 36001 63532
rect 36035 63529 36047 63563
rect 35989 63523 36047 63529
rect 36078 63520 36084 63572
rect 36136 63560 36142 63572
rect 36630 63560 36636 63572
rect 36136 63532 36636 63560
rect 36136 63520 36142 63532
rect 36630 63520 36636 63532
rect 36688 63560 36694 63572
rect 36725 63563 36783 63569
rect 36725 63560 36737 63563
rect 36688 63532 36737 63560
rect 36688 63520 36694 63532
rect 36725 63529 36737 63532
rect 36771 63529 36783 63563
rect 36725 63523 36783 63529
rect 25314 63452 25320 63504
rect 25372 63492 25378 63504
rect 61562 63492 61568 63504
rect 25372 63464 61568 63492
rect 25372 63452 25378 63464
rect 61562 63452 61568 63464
rect 61620 63452 61626 63504
rect 35342 63384 35348 63436
rect 35400 63424 35406 63436
rect 36446 63424 36452 63436
rect 35400 63396 36452 63424
rect 35400 63384 35406 63396
rect 36446 63384 36452 63396
rect 36504 63384 36510 63436
rect 37001 63427 37059 63433
rect 37001 63393 37013 63427
rect 37047 63424 37059 63427
rect 37274 63424 37280 63436
rect 37047 63396 37280 63424
rect 37047 63393 37059 63396
rect 37001 63387 37059 63393
rect 37274 63384 37280 63396
rect 37332 63424 37338 63436
rect 38010 63424 38016 63436
rect 37332 63396 38016 63424
rect 37332 63384 37338 63396
rect 38010 63384 38016 63396
rect 38068 63384 38074 63436
rect 66254 63424 66260 63436
rect 66215 63396 66260 63424
rect 66254 63384 66260 63396
rect 66312 63384 66318 63436
rect 1394 63356 1400 63368
rect 1355 63328 1400 63356
rect 1394 63316 1400 63328
rect 1452 63316 1458 63368
rect 24394 63316 24400 63368
rect 24452 63356 24458 63368
rect 24489 63359 24547 63365
rect 24489 63356 24501 63359
rect 24452 63328 24501 63356
rect 24452 63316 24458 63328
rect 24489 63325 24501 63328
rect 24535 63325 24547 63359
rect 24489 63319 24547 63325
rect 34885 63359 34943 63365
rect 34885 63325 34897 63359
rect 34931 63325 34943 63359
rect 34885 63319 34943 63325
rect 35621 63359 35679 63365
rect 35621 63325 35633 63359
rect 35667 63356 35679 63359
rect 35710 63356 35716 63368
rect 35667 63328 35716 63356
rect 35667 63325 35679 63328
rect 35621 63319 35679 63325
rect 1673 63291 1731 63297
rect 1673 63257 1685 63291
rect 1719 63288 1731 63291
rect 24854 63288 24860 63300
rect 1719 63260 6914 63288
rect 24815 63260 24860 63288
rect 1719 63257 1731 63260
rect 1673 63251 1731 63257
rect 6886 63220 6914 63260
rect 24854 63248 24860 63260
rect 24912 63248 24918 63300
rect 34900 63288 34928 63319
rect 35710 63316 35716 63328
rect 35768 63316 35774 63368
rect 36814 63316 36820 63368
rect 36872 63356 36878 63368
rect 36909 63359 36967 63365
rect 36909 63356 36921 63359
rect 36872 63328 36921 63356
rect 36872 63316 36878 63328
rect 36909 63325 36921 63328
rect 36955 63325 36967 63359
rect 36909 63319 36967 63325
rect 37093 63359 37151 63365
rect 37093 63325 37105 63359
rect 37139 63325 37151 63359
rect 37093 63319 37151 63325
rect 37185 63359 37243 63365
rect 37185 63325 37197 63359
rect 37231 63356 37243 63359
rect 37734 63356 37740 63368
rect 37231 63328 37740 63356
rect 37231 63325 37243 63328
rect 37185 63319 37243 63325
rect 34900 63260 36216 63288
rect 31938 63220 31944 63232
rect 6886 63192 31944 63220
rect 31938 63180 31944 63192
rect 31996 63180 32002 63232
rect 35989 63223 36047 63229
rect 35989 63189 36001 63223
rect 36035 63220 36047 63223
rect 36078 63220 36084 63232
rect 36035 63192 36084 63220
rect 36035 63189 36047 63192
rect 35989 63183 36047 63189
rect 36078 63180 36084 63192
rect 36136 63180 36142 63232
rect 36188 63229 36216 63260
rect 36630 63248 36636 63300
rect 36688 63288 36694 63300
rect 37108 63288 37136 63319
rect 37734 63316 37740 63328
rect 37792 63316 37798 63368
rect 68094 63356 68100 63368
rect 68055 63328 68100 63356
rect 68094 63316 68100 63328
rect 68152 63316 68158 63368
rect 66438 63288 66444 63300
rect 36688 63260 37136 63288
rect 66399 63260 66444 63288
rect 36688 63248 36694 63260
rect 66438 63248 66444 63260
rect 66496 63248 66502 63300
rect 36173 63223 36231 63229
rect 36173 63189 36185 63223
rect 36219 63189 36231 63223
rect 36173 63183 36231 63189
rect 1104 63130 68816 63152
rect 1104 63078 19574 63130
rect 19626 63078 19638 63130
rect 19690 63078 19702 63130
rect 19754 63078 19766 63130
rect 19818 63078 19830 63130
rect 19882 63078 50294 63130
rect 50346 63078 50358 63130
rect 50410 63078 50422 63130
rect 50474 63078 50486 63130
rect 50538 63078 50550 63130
rect 50602 63078 68816 63130
rect 1104 63056 68816 63078
rect 56226 63016 56232 63028
rect 24504 62988 56232 63016
rect 23106 62880 23112 62892
rect 23019 62852 23112 62880
rect 23106 62840 23112 62852
rect 23164 62880 23170 62892
rect 23382 62880 23388 62892
rect 23164 62852 23388 62880
rect 23164 62840 23170 62852
rect 23382 62840 23388 62852
rect 23440 62840 23446 62892
rect 23477 62883 23535 62889
rect 23477 62849 23489 62883
rect 23523 62880 23535 62883
rect 24121 62883 24179 62889
rect 24121 62880 24133 62883
rect 23523 62852 24133 62880
rect 23523 62849 23535 62852
rect 23477 62843 23535 62849
rect 24121 62849 24133 62852
rect 24167 62880 24179 62883
rect 24394 62880 24400 62892
rect 24167 62852 24400 62880
rect 24167 62849 24179 62852
rect 24121 62843 24179 62849
rect 24394 62840 24400 62852
rect 24452 62840 24458 62892
rect 23842 62772 23848 62824
rect 23900 62812 23906 62824
rect 24504 62821 24532 62988
rect 56226 62976 56232 62988
rect 56284 62976 56290 63028
rect 66438 62976 66444 63028
rect 66496 63016 66502 63028
rect 67545 63019 67603 63025
rect 67545 63016 67557 63019
rect 66496 62988 67557 63016
rect 66496 62976 66502 62988
rect 67545 62985 67557 62988
rect 67591 62985 67603 63019
rect 67545 62979 67603 62985
rect 24854 62908 24860 62960
rect 24912 62948 24918 62960
rect 28537 62951 28595 62957
rect 24912 62920 28488 62948
rect 24912 62908 24918 62920
rect 28460 62889 28488 62920
rect 28537 62917 28549 62951
rect 28583 62948 28595 62951
rect 29273 62951 29331 62957
rect 29273 62948 29285 62951
rect 28583 62920 29285 62948
rect 28583 62917 28595 62920
rect 28537 62911 28595 62917
rect 29273 62917 29285 62920
rect 29319 62917 29331 62951
rect 35342 62948 35348 62960
rect 35303 62920 35348 62948
rect 29273 62911 29331 62917
rect 35342 62908 35348 62920
rect 35400 62908 35406 62960
rect 35434 62908 35440 62960
rect 35492 62948 35498 62960
rect 35545 62951 35603 62957
rect 35545 62948 35557 62951
rect 35492 62920 35557 62948
rect 35492 62908 35498 62920
rect 35545 62917 35557 62920
rect 35591 62917 35603 62951
rect 44174 62948 44180 62960
rect 35545 62911 35603 62917
rect 35866 62920 44180 62948
rect 28445 62883 28503 62889
rect 28445 62849 28457 62883
rect 28491 62849 28503 62883
rect 28445 62843 28503 62849
rect 34793 62883 34851 62889
rect 34793 62849 34805 62883
rect 34839 62880 34851 62883
rect 35866 62880 35894 62920
rect 44174 62908 44180 62920
rect 44232 62908 44238 62960
rect 34839 62852 35894 62880
rect 36173 62883 36231 62889
rect 34839 62849 34851 62852
rect 34793 62843 34851 62849
rect 36173 62849 36185 62883
rect 36219 62880 36231 62883
rect 36354 62880 36360 62892
rect 36219 62852 36360 62880
rect 36219 62849 36231 62852
rect 36173 62843 36231 62849
rect 24489 62815 24547 62821
rect 24489 62812 24501 62815
rect 23900 62784 24501 62812
rect 23900 62772 23906 62784
rect 24489 62781 24501 62784
rect 24535 62781 24547 62815
rect 24489 62775 24547 62781
rect 28460 62744 28488 62843
rect 36354 62840 36360 62852
rect 36412 62840 36418 62892
rect 36446 62840 36452 62892
rect 36504 62880 36510 62892
rect 37642 62880 37648 62892
rect 36504 62852 36549 62880
rect 37603 62852 37648 62880
rect 36504 62840 36510 62852
rect 37642 62840 37648 62852
rect 37700 62840 37706 62892
rect 37829 62883 37887 62889
rect 37829 62849 37841 62883
rect 37875 62849 37887 62883
rect 37829 62843 37887 62849
rect 29086 62812 29092 62824
rect 29047 62784 29092 62812
rect 29086 62772 29092 62784
rect 29144 62772 29150 62824
rect 29270 62772 29276 62824
rect 29328 62812 29334 62824
rect 29549 62815 29607 62821
rect 29549 62812 29561 62815
rect 29328 62784 29561 62812
rect 29328 62772 29334 62784
rect 29549 62781 29561 62784
rect 29595 62781 29607 62815
rect 32950 62812 32956 62824
rect 32911 62784 32956 62812
rect 29549 62775 29607 62781
rect 32950 62772 32956 62784
rect 33008 62772 33014 62824
rect 33134 62812 33140 62824
rect 33095 62784 33140 62812
rect 33134 62772 33140 62784
rect 33192 62772 33198 62824
rect 36078 62812 36084 62824
rect 35544 62784 36084 62812
rect 32490 62744 32496 62756
rect 28460 62716 32496 62744
rect 32490 62704 32496 62716
rect 32548 62704 32554 62756
rect 35434 62636 35440 62688
rect 35492 62676 35498 62688
rect 35544 62685 35572 62784
rect 36078 62772 36084 62784
rect 36136 62772 36142 62824
rect 36262 62812 36268 62824
rect 36223 62784 36268 62812
rect 36262 62772 36268 62784
rect 36320 62772 36326 62824
rect 35710 62744 35716 62756
rect 35671 62716 35716 62744
rect 35710 62704 35716 62716
rect 35768 62744 35774 62756
rect 36630 62744 36636 62756
rect 35768 62716 35894 62744
rect 36591 62716 36636 62744
rect 35768 62704 35774 62716
rect 35529 62679 35587 62685
rect 35529 62676 35541 62679
rect 35492 62648 35541 62676
rect 35492 62636 35498 62648
rect 35529 62645 35541 62648
rect 35575 62645 35587 62679
rect 35866 62676 35894 62716
rect 36630 62704 36636 62716
rect 36688 62704 36694 62756
rect 37844 62744 37872 62843
rect 37918 62840 37924 62892
rect 37976 62880 37982 62892
rect 38545 62883 38603 62889
rect 38545 62880 38557 62883
rect 37976 62852 38557 62880
rect 37976 62840 37982 62852
rect 38545 62849 38557 62852
rect 38591 62849 38603 62883
rect 38545 62843 38603 62849
rect 57238 62840 57244 62892
rect 57296 62880 57302 62892
rect 67453 62883 67511 62889
rect 67453 62880 67465 62883
rect 57296 62852 67465 62880
rect 57296 62840 57302 62852
rect 67453 62849 67465 62852
rect 67499 62880 67511 62883
rect 67542 62880 67548 62892
rect 67499 62852 67548 62880
rect 67499 62849 67511 62852
rect 67453 62843 67511 62849
rect 67542 62840 67548 62852
rect 67600 62840 67606 62892
rect 38102 62772 38108 62824
rect 38160 62812 38166 62824
rect 38289 62815 38347 62821
rect 38289 62812 38301 62815
rect 38160 62784 38301 62812
rect 38160 62772 38166 62784
rect 38289 62781 38301 62784
rect 38335 62781 38347 62815
rect 38289 62775 38347 62781
rect 38010 62744 38016 62756
rect 37844 62716 38016 62744
rect 38010 62704 38016 62716
rect 38068 62744 38074 62756
rect 38068 62716 38332 62744
rect 38068 62704 38074 62716
rect 35986 62676 35992 62688
rect 35866 62648 35992 62676
rect 35529 62639 35587 62645
rect 35986 62636 35992 62648
rect 36044 62636 36050 62688
rect 36170 62636 36176 62688
rect 36228 62676 36234 62688
rect 37737 62679 37795 62685
rect 36228 62648 36273 62676
rect 36228 62636 36234 62648
rect 37737 62645 37749 62679
rect 37783 62676 37795 62679
rect 38194 62676 38200 62688
rect 37783 62648 38200 62676
rect 37783 62645 37795 62648
rect 37737 62639 37795 62645
rect 38194 62636 38200 62648
rect 38252 62636 38258 62688
rect 38304 62676 38332 62716
rect 39669 62679 39727 62685
rect 39669 62676 39681 62679
rect 38304 62648 39681 62676
rect 39669 62645 39681 62648
rect 39715 62645 39727 62679
rect 39669 62639 39727 62645
rect 1104 62586 68816 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 34934 62586
rect 34986 62534 34998 62586
rect 35050 62534 35062 62586
rect 35114 62534 35126 62586
rect 35178 62534 35190 62586
rect 35242 62534 65654 62586
rect 65706 62534 65718 62586
rect 65770 62534 65782 62586
rect 65834 62534 65846 62586
rect 65898 62534 65910 62586
rect 65962 62534 68816 62586
rect 1104 62512 68816 62534
rect 23106 62432 23112 62484
rect 23164 62472 23170 62484
rect 31018 62472 31024 62484
rect 23164 62444 31024 62472
rect 23164 62432 23170 62444
rect 31018 62432 31024 62444
rect 31076 62432 31082 62484
rect 33134 62472 33140 62484
rect 33095 62444 33140 62472
rect 33134 62432 33140 62444
rect 33192 62432 33198 62484
rect 37737 62475 37795 62481
rect 37737 62441 37749 62475
rect 37783 62472 37795 62475
rect 37918 62472 37924 62484
rect 37783 62444 37924 62472
rect 37783 62441 37795 62444
rect 37737 62435 37795 62441
rect 37918 62432 37924 62444
rect 37976 62432 37982 62484
rect 35986 62364 35992 62416
rect 36044 62404 36050 62416
rect 37642 62404 37648 62416
rect 36044 62376 37648 62404
rect 36044 62364 36050 62376
rect 37642 62364 37648 62376
rect 37700 62404 37706 62416
rect 37700 62376 38148 62404
rect 37700 62364 37706 62376
rect 23106 62336 23112 62348
rect 23067 62308 23112 62336
rect 23106 62296 23112 62308
rect 23164 62296 23170 62348
rect 29362 62296 29368 62348
rect 29420 62336 29426 62348
rect 30837 62339 30895 62345
rect 30837 62336 30849 62339
rect 29420 62308 30849 62336
rect 29420 62296 29426 62308
rect 30837 62305 30849 62308
rect 30883 62305 30895 62339
rect 35434 62336 35440 62348
rect 30837 62299 30895 62305
rect 35268 62308 35440 62336
rect 19889 62271 19947 62277
rect 19889 62237 19901 62271
rect 19935 62268 19947 62271
rect 21818 62268 21824 62280
rect 19935 62240 21824 62268
rect 19935 62237 19947 62240
rect 19889 62231 19947 62237
rect 21818 62228 21824 62240
rect 21876 62228 21882 62280
rect 22649 62271 22707 62277
rect 22649 62237 22661 62271
rect 22695 62268 22707 62271
rect 24394 62268 24400 62280
rect 22695 62240 24400 62268
rect 22695 62237 22707 62240
rect 22649 62231 22707 62237
rect 24394 62228 24400 62240
rect 24452 62228 24458 62280
rect 26234 62228 26240 62280
rect 26292 62268 26298 62280
rect 28077 62271 28135 62277
rect 28077 62268 28089 62271
rect 26292 62240 26337 62268
rect 26436 62240 28089 62268
rect 26292 62228 26298 62240
rect 25314 62200 25320 62212
rect 25275 62172 25320 62200
rect 25314 62160 25320 62172
rect 25372 62160 25378 62212
rect 25958 62160 25964 62212
rect 26016 62200 26022 62212
rect 26436 62200 26464 62240
rect 28077 62237 28089 62240
rect 28123 62237 28135 62271
rect 28994 62268 29000 62280
rect 28955 62240 29000 62268
rect 28077 62231 28135 62237
rect 28994 62228 29000 62240
rect 29052 62228 29058 62280
rect 29730 62268 29736 62280
rect 29691 62240 29736 62268
rect 29730 62228 29736 62240
rect 29788 62228 29794 62280
rect 30374 62268 30380 62280
rect 30335 62240 30380 62268
rect 30374 62228 30380 62240
rect 30432 62228 30438 62280
rect 33045 62271 33103 62277
rect 33045 62237 33057 62271
rect 33091 62237 33103 62271
rect 33045 62231 33103 62237
rect 26510 62209 26516 62212
rect 26016 62172 26464 62200
rect 26016 62160 26022 62172
rect 26504 62163 26516 62209
rect 26568 62200 26574 62212
rect 29825 62203 29883 62209
rect 26568 62172 26604 62200
rect 26510 62160 26516 62163
rect 26568 62160 26574 62172
rect 29825 62169 29837 62203
rect 29871 62200 29883 62203
rect 30561 62203 30619 62209
rect 30561 62200 30573 62203
rect 29871 62172 30573 62200
rect 29871 62169 29883 62172
rect 29825 62163 29883 62169
rect 30561 62169 30573 62172
rect 30607 62169 30619 62203
rect 30561 62163 30619 62169
rect 19334 62092 19340 62144
rect 19392 62132 19398 62144
rect 19889 62135 19947 62141
rect 19889 62132 19901 62135
rect 19392 62104 19901 62132
rect 19392 62092 19398 62104
rect 19889 62101 19901 62104
rect 19935 62101 19947 62135
rect 19889 62095 19947 62101
rect 27430 62092 27436 62144
rect 27488 62132 27494 62144
rect 27617 62135 27675 62141
rect 27617 62132 27629 62135
rect 27488 62104 27629 62132
rect 27488 62092 27494 62104
rect 27617 62101 27629 62104
rect 27663 62101 27675 62135
rect 28258 62132 28264 62144
rect 28219 62104 28264 62132
rect 27617 62095 27675 62101
rect 28258 62092 28264 62104
rect 28316 62092 28322 62144
rect 28810 62132 28816 62144
rect 28771 62104 28816 62132
rect 28810 62092 28816 62104
rect 28868 62092 28874 62144
rect 29730 62092 29736 62144
rect 29788 62132 29794 62144
rect 33060 62132 33088 62231
rect 34698 62228 34704 62280
rect 34756 62268 34762 62280
rect 35268 62277 35296 62308
rect 35434 62296 35440 62308
rect 35492 62296 35498 62348
rect 35529 62339 35587 62345
rect 35529 62305 35541 62339
rect 35575 62336 35587 62339
rect 36630 62336 36636 62348
rect 35575 62308 36636 62336
rect 35575 62305 35587 62308
rect 35529 62299 35587 62305
rect 36630 62296 36636 62308
rect 36688 62296 36694 62348
rect 35253 62271 35311 62277
rect 35253 62268 35265 62271
rect 34756 62240 35265 62268
rect 34756 62228 34762 62240
rect 35253 62237 35265 62240
rect 35299 62237 35311 62271
rect 35253 62231 35311 62237
rect 35342 62228 35348 62280
rect 35400 62268 35406 62280
rect 38010 62268 38016 62280
rect 35400 62240 35445 62268
rect 37971 62240 38016 62268
rect 35400 62228 35406 62240
rect 38010 62228 38016 62240
rect 38068 62228 38074 62280
rect 38120 62277 38148 62376
rect 38105 62271 38163 62277
rect 38105 62237 38117 62271
rect 38151 62237 38163 62271
rect 38105 62231 38163 62237
rect 38194 62228 38200 62280
rect 38252 62268 38258 62280
rect 38381 62271 38439 62277
rect 38252 62240 38297 62268
rect 38252 62228 38258 62240
rect 38381 62237 38393 62271
rect 38427 62237 38439 62271
rect 38381 62231 38439 62237
rect 36630 62160 36636 62212
rect 36688 62200 36694 62212
rect 38396 62200 38424 62231
rect 66254 62228 66260 62280
rect 66312 62268 66318 62280
rect 67913 62271 67971 62277
rect 67913 62268 67925 62271
rect 66312 62240 67925 62268
rect 66312 62228 66318 62240
rect 67913 62237 67925 62240
rect 67959 62237 67971 62271
rect 67913 62231 67971 62237
rect 36688 62172 38424 62200
rect 36688 62160 36694 62172
rect 33686 62132 33692 62144
rect 29788 62104 33692 62132
rect 29788 62092 29794 62104
rect 33686 62092 33692 62104
rect 33744 62092 33750 62144
rect 35526 62132 35532 62144
rect 35487 62104 35532 62132
rect 35526 62092 35532 62104
rect 35584 62092 35590 62144
rect 1104 62042 68816 62064
rect 1104 61990 19574 62042
rect 19626 61990 19638 62042
rect 19690 61990 19702 62042
rect 19754 61990 19766 62042
rect 19818 61990 19830 62042
rect 19882 61990 50294 62042
rect 50346 61990 50358 62042
rect 50410 61990 50422 62042
rect 50474 61990 50486 62042
rect 50538 61990 50550 62042
rect 50602 61990 68816 62042
rect 1104 61968 68816 61990
rect 19334 61888 19340 61940
rect 19392 61888 19398 61940
rect 26145 61931 26203 61937
rect 26145 61897 26157 61931
rect 26191 61928 26203 61931
rect 26234 61928 26240 61940
rect 26191 61900 26240 61928
rect 26191 61897 26203 61900
rect 26145 61891 26203 61897
rect 26234 61888 26240 61900
rect 26292 61888 26298 61940
rect 38930 61928 38936 61940
rect 27448 61900 38936 61928
rect 2958 61820 2964 61872
rect 3016 61860 3022 61872
rect 19352 61860 19380 61888
rect 25130 61860 25136 61872
rect 3016 61832 6914 61860
rect 3016 61820 3022 61832
rect 6886 61588 6914 61832
rect 19260 61832 19380 61860
rect 22066 61832 24256 61860
rect 25043 61832 25136 61860
rect 19260 61801 19288 61832
rect 19245 61795 19303 61801
rect 19245 61761 19257 61795
rect 19291 61761 19303 61795
rect 19245 61755 19303 61761
rect 19334 61752 19340 61804
rect 19392 61792 19398 61804
rect 19501 61795 19559 61801
rect 19501 61792 19513 61795
rect 19392 61764 19513 61792
rect 19392 61752 19398 61764
rect 19501 61761 19513 61764
rect 19547 61761 19559 61795
rect 19501 61755 19559 61761
rect 20714 61752 20720 61804
rect 20772 61792 20778 61804
rect 21269 61795 21327 61801
rect 21269 61792 21281 61795
rect 20772 61764 21281 61792
rect 20772 61752 20778 61764
rect 21269 61761 21281 61764
rect 21315 61761 21327 61795
rect 21818 61792 21824 61804
rect 21779 61764 21824 61792
rect 21269 61755 21327 61761
rect 21818 61752 21824 61764
rect 21876 61792 21882 61804
rect 22066 61792 22094 61832
rect 21876 61764 22094 61792
rect 24228 61792 24256 61832
rect 25130 61820 25136 61832
rect 25188 61860 25194 61872
rect 26050 61860 26056 61872
rect 25188 61832 26056 61860
rect 25188 61820 25194 61832
rect 26050 61820 26056 61832
rect 26108 61820 26114 61872
rect 25682 61792 25688 61804
rect 24228 61764 25688 61792
rect 21876 61752 21882 61764
rect 25682 61752 25688 61764
rect 25740 61792 25746 61804
rect 25958 61792 25964 61804
rect 25740 61764 25964 61792
rect 25740 61752 25746 61764
rect 25958 61752 25964 61764
rect 26016 61752 26022 61804
rect 22738 61724 22744 61736
rect 22699 61696 22744 61724
rect 22738 61684 22744 61696
rect 22796 61684 22802 61736
rect 22925 61727 22983 61733
rect 22925 61693 22937 61727
rect 22971 61724 22983 61727
rect 23566 61724 23572 61736
rect 22971 61696 23572 61724
rect 22971 61693 22983 61696
rect 22925 61687 22983 61693
rect 23566 61684 23572 61696
rect 23624 61684 23630 61736
rect 23661 61727 23719 61733
rect 23661 61693 23673 61727
rect 23707 61693 23719 61727
rect 23661 61687 23719 61693
rect 23676 61656 23704 61687
rect 25866 61684 25872 61736
rect 25924 61724 25930 61736
rect 27448 61724 27476 61900
rect 38930 61888 38936 61900
rect 38988 61888 38994 61940
rect 27792 61863 27850 61869
rect 27792 61829 27804 61863
rect 27838 61860 27850 61863
rect 28810 61860 28816 61872
rect 27838 61832 28816 61860
rect 27838 61829 27850 61832
rect 27792 61823 27850 61829
rect 28810 61820 28816 61832
rect 28868 61820 28874 61872
rect 31754 61860 31760 61872
rect 29656 61832 31760 61860
rect 27525 61795 27583 61801
rect 27525 61761 27537 61795
rect 27571 61792 27583 61795
rect 28258 61792 28264 61804
rect 27571 61764 28264 61792
rect 27571 61761 27583 61764
rect 27525 61755 27583 61761
rect 28258 61752 28264 61764
rect 28316 61752 28322 61804
rect 29656 61801 29684 61832
rect 31754 61820 31760 61832
rect 31812 61820 31818 61872
rect 66254 61860 66260 61872
rect 65812 61832 66260 61860
rect 29641 61795 29699 61801
rect 29641 61761 29653 61795
rect 29687 61761 29699 61795
rect 29641 61755 29699 61761
rect 29908 61795 29966 61801
rect 29908 61761 29920 61795
rect 29954 61792 29966 61795
rect 30282 61792 30288 61804
rect 29954 61764 30288 61792
rect 29954 61761 29966 61764
rect 29908 61755 29966 61761
rect 30282 61752 30288 61764
rect 30340 61752 30346 61804
rect 33680 61795 33738 61801
rect 33680 61761 33692 61795
rect 33726 61792 33738 61795
rect 34790 61792 34796 61804
rect 33726 61764 34796 61792
rect 33726 61761 33738 61764
rect 33680 61755 33738 61761
rect 34790 61752 34796 61764
rect 34848 61752 34854 61804
rect 35989 61795 36047 61801
rect 35989 61792 36001 61795
rect 35360 61764 36001 61792
rect 33410 61724 33416 61736
rect 25924 61696 27476 61724
rect 33371 61696 33416 61724
rect 25924 61684 25930 61696
rect 33410 61684 33416 61696
rect 33468 61684 33474 61736
rect 35360 61724 35388 61764
rect 35989 61761 36001 61764
rect 36035 61761 36047 61795
rect 35989 61755 36047 61761
rect 36265 61795 36323 61801
rect 36265 61761 36277 61795
rect 36311 61792 36323 61795
rect 36446 61792 36452 61804
rect 36311 61764 36452 61792
rect 36311 61761 36323 61764
rect 36265 61755 36323 61761
rect 36446 61752 36452 61764
rect 36504 61752 36510 61804
rect 65812 61801 65840 61832
rect 66254 61820 66260 61832
rect 66312 61820 66318 61872
rect 67634 61860 67640 61872
rect 67595 61832 67640 61860
rect 67634 61820 67640 61832
rect 67692 61820 67698 61872
rect 65797 61795 65855 61801
rect 65797 61761 65809 61795
rect 65843 61761 65855 61795
rect 65797 61755 65855 61761
rect 35802 61724 35808 61736
rect 34808 61696 35388 61724
rect 35763 61696 35808 61724
rect 20180 61628 23704 61656
rect 20180 61588 20208 61628
rect 6886 61560 20208 61588
rect 20346 61548 20352 61600
rect 20404 61588 20410 61600
rect 20625 61591 20683 61597
rect 20625 61588 20637 61591
rect 20404 61560 20637 61588
rect 20404 61548 20410 61560
rect 20625 61557 20637 61560
rect 20671 61557 20683 61591
rect 21082 61588 21088 61600
rect 21043 61560 21088 61588
rect 20625 61551 20683 61557
rect 21082 61548 21088 61560
rect 21140 61548 21146 61600
rect 21174 61548 21180 61600
rect 21232 61588 21238 61600
rect 21821 61591 21879 61597
rect 21821 61588 21833 61591
rect 21232 61560 21833 61588
rect 21232 61548 21238 61560
rect 21821 61557 21833 61560
rect 21867 61557 21879 61591
rect 21821 61551 21879 61557
rect 24302 61548 24308 61600
rect 24360 61588 24366 61600
rect 25225 61591 25283 61597
rect 25225 61588 25237 61591
rect 24360 61560 25237 61588
rect 24360 61548 24366 61560
rect 25225 61557 25237 61560
rect 25271 61588 25283 61591
rect 27798 61588 27804 61600
rect 25271 61560 27804 61588
rect 25271 61557 25283 61560
rect 25225 61551 25283 61557
rect 27798 61548 27804 61560
rect 27856 61548 27862 61600
rect 27890 61548 27896 61600
rect 27948 61588 27954 61600
rect 28905 61591 28963 61597
rect 28905 61588 28917 61591
rect 27948 61560 28917 61588
rect 27948 61548 27954 61560
rect 28905 61557 28917 61560
rect 28951 61557 28963 61591
rect 28905 61551 28963 61557
rect 30374 61548 30380 61600
rect 30432 61588 30438 61600
rect 31021 61591 31079 61597
rect 31021 61588 31033 61591
rect 30432 61560 31033 61588
rect 30432 61548 30438 61560
rect 31021 61557 31033 61560
rect 31067 61557 31079 61591
rect 31021 61551 31079 61557
rect 34698 61548 34704 61600
rect 34756 61588 34762 61600
rect 34808 61597 34836 61696
rect 35802 61684 35808 61696
rect 35860 61684 35866 61736
rect 36078 61724 36084 61736
rect 36039 61696 36084 61724
rect 36078 61684 36084 61696
rect 36136 61684 36142 61736
rect 36173 61727 36231 61733
rect 36173 61693 36185 61727
rect 36219 61693 36231 61727
rect 36173 61687 36231 61693
rect 65981 61727 66039 61733
rect 65981 61693 65993 61727
rect 66027 61724 66039 61727
rect 67634 61724 67640 61736
rect 66027 61696 67640 61724
rect 66027 61693 66039 61696
rect 65981 61687 66039 61693
rect 35986 61616 35992 61668
rect 36044 61656 36050 61668
rect 36188 61656 36216 61687
rect 67634 61684 67640 61696
rect 67692 61684 67698 61736
rect 36044 61628 36216 61656
rect 36044 61616 36050 61628
rect 34793 61591 34851 61597
rect 34793 61588 34805 61591
rect 34756 61560 34805 61588
rect 34756 61548 34762 61560
rect 34793 61557 34805 61560
rect 34839 61557 34851 61591
rect 34793 61551 34851 61557
rect 1104 61498 68816 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 34934 61498
rect 34986 61446 34998 61498
rect 35050 61446 35062 61498
rect 35114 61446 35126 61498
rect 35178 61446 35190 61498
rect 35242 61446 65654 61498
rect 65706 61446 65718 61498
rect 65770 61446 65782 61498
rect 65834 61446 65846 61498
rect 65898 61446 65910 61498
rect 65962 61446 68816 61498
rect 1104 61424 68816 61446
rect 20346 61384 20352 61396
rect 19444 61356 20352 61384
rect 19444 61260 19472 61356
rect 20346 61344 20352 61356
rect 20404 61344 20410 61396
rect 20714 61384 20720 61396
rect 20675 61356 20720 61384
rect 20714 61344 20720 61356
rect 20772 61344 20778 61396
rect 23566 61384 23572 61396
rect 23527 61356 23572 61384
rect 23566 61344 23572 61356
rect 23624 61344 23630 61396
rect 26421 61387 26479 61393
rect 26421 61353 26433 61387
rect 26467 61384 26479 61387
rect 26510 61384 26516 61396
rect 26467 61356 26516 61384
rect 26467 61353 26479 61356
rect 26421 61347 26479 61353
rect 26510 61344 26516 61356
rect 26568 61344 26574 61396
rect 28629 61387 28687 61393
rect 28629 61353 28641 61387
rect 28675 61384 28687 61387
rect 28994 61384 29000 61396
rect 28675 61356 29000 61384
rect 28675 61353 28687 61356
rect 28629 61347 28687 61353
rect 28994 61344 29000 61356
rect 29052 61344 29058 61396
rect 32950 61384 32956 61396
rect 30852 61356 32956 61384
rect 19610 61276 19616 61328
rect 19668 61316 19674 61328
rect 19668 61288 20760 61316
rect 19668 61276 19674 61288
rect 19426 61248 19432 61260
rect 19339 61220 19432 61248
rect 19426 61208 19432 61220
rect 19484 61208 19490 61260
rect 20349 61251 20407 61257
rect 20349 61217 20361 61251
rect 20395 61217 20407 61251
rect 20349 61211 20407 61217
rect 18230 61140 18236 61192
rect 18288 61180 18294 61192
rect 19610 61180 19616 61192
rect 18288 61152 19616 61180
rect 18288 61140 18294 61152
rect 19610 61140 19616 61152
rect 19668 61140 19674 61192
rect 20364 61182 20392 61211
rect 20272 61154 20392 61182
rect 20533 61183 20591 61189
rect 19797 61047 19855 61053
rect 19797 61013 19809 61047
rect 19843 61044 19855 61047
rect 19978 61044 19984 61056
rect 19843 61016 19984 61044
rect 19843 61013 19855 61016
rect 19797 61007 19855 61013
rect 19978 61004 19984 61016
rect 20036 61004 20042 61056
rect 20272 61044 20300 61154
rect 20533 61149 20545 61183
rect 20579 61180 20591 61183
rect 20732 61180 20760 61288
rect 27798 61276 27804 61328
rect 27856 61316 27862 61328
rect 29730 61316 29736 61328
rect 27856 61288 29736 61316
rect 27856 61276 27862 61288
rect 29730 61276 29736 61288
rect 29788 61276 29794 61328
rect 21174 61248 21180 61260
rect 21135 61220 21180 61248
rect 21174 61208 21180 61220
rect 21232 61208 21238 61260
rect 24854 61248 24860 61260
rect 23492 61220 24860 61248
rect 20579 61152 20760 61180
rect 20579 61149 20591 61152
rect 20533 61143 20591 61149
rect 21082 61140 21088 61192
rect 21140 61180 21146 61192
rect 23492 61189 23520 61220
rect 24854 61208 24860 61220
rect 24912 61208 24918 61260
rect 27709 61251 27767 61257
rect 27709 61248 27721 61251
rect 26620 61220 27721 61248
rect 21433 61183 21491 61189
rect 21433 61180 21445 61183
rect 21140 61152 21445 61180
rect 21140 61140 21146 61152
rect 21433 61149 21445 61152
rect 21479 61149 21491 61183
rect 21433 61143 21491 61149
rect 23477 61183 23535 61189
rect 23477 61149 23489 61183
rect 23523 61149 23535 61183
rect 24394 61180 24400 61192
rect 24355 61152 24400 61180
rect 23477 61143 23535 61149
rect 24394 61140 24400 61152
rect 24452 61140 24458 61192
rect 26620 61189 26648 61220
rect 27709 61217 27721 61220
rect 27755 61217 27767 61251
rect 27709 61211 27767 61217
rect 26605 61183 26663 61189
rect 26605 61149 26617 61183
rect 26651 61149 26663 61183
rect 27430 61180 27436 61192
rect 27391 61152 27436 61180
rect 26605 61143 26663 61149
rect 27430 61140 27436 61152
rect 27488 61140 27494 61192
rect 27525 61183 27583 61189
rect 27525 61149 27537 61183
rect 27571 61149 27583 61183
rect 27525 61143 27583 61149
rect 25225 61115 25283 61121
rect 25225 61081 25237 61115
rect 25271 61112 25283 61115
rect 25866 61112 25872 61124
rect 25271 61084 25872 61112
rect 25271 61081 25283 61084
rect 25225 61075 25283 61081
rect 25866 61072 25872 61084
rect 25924 61072 25930 61124
rect 27540 61112 27568 61143
rect 27890 61140 27896 61192
rect 27948 61180 27954 61192
rect 28261 61183 28319 61189
rect 28261 61180 28273 61183
rect 27948 61152 28273 61180
rect 27948 61140 27954 61152
rect 28261 61149 28273 61152
rect 28307 61149 28319 61183
rect 28261 61143 28319 61149
rect 28350 61140 28356 61192
rect 28408 61180 28414 61192
rect 30852 61189 30880 61356
rect 32950 61344 32956 61356
rect 33008 61384 33014 61396
rect 33045 61387 33103 61393
rect 33045 61384 33057 61387
rect 33008 61356 33057 61384
rect 33008 61344 33014 61356
rect 33045 61353 33057 61356
rect 33091 61353 33103 61387
rect 33045 61347 33103 61353
rect 33410 61344 33416 61396
rect 33468 61384 33474 61396
rect 67634 61384 67640 61396
rect 33468 61356 36860 61384
rect 67595 61356 67640 61384
rect 33468 61344 33474 61356
rect 34790 61316 34796 61328
rect 34751 61288 34796 61316
rect 34790 61276 34796 61288
rect 34848 61276 34854 61328
rect 36078 61276 36084 61328
rect 36136 61276 36142 61328
rect 31478 61248 31484 61260
rect 30944 61220 31484 61248
rect 30944 61189 30972 61220
rect 31478 61208 31484 61220
rect 31536 61208 31542 61260
rect 28445 61183 28503 61189
rect 28445 61180 28457 61183
rect 28408 61152 28457 61180
rect 28408 61140 28414 61152
rect 28445 61149 28457 61152
rect 28491 61149 28503 61183
rect 28445 61143 28503 61149
rect 30817 61183 30880 61189
rect 30817 61149 30829 61183
rect 30863 61152 30880 61183
rect 30910 61183 30972 61189
rect 30863 61149 30875 61152
rect 30817 61143 30875 61149
rect 30910 61149 30922 61183
rect 30956 61152 30972 61183
rect 30956 61149 30968 61152
rect 30910 61143 30968 61149
rect 31018 61140 31024 61192
rect 31076 61180 31082 61192
rect 31076 61152 31121 61180
rect 31076 61140 31082 61152
rect 31202 61140 31208 61192
rect 31260 61180 31266 61192
rect 31665 61183 31723 61189
rect 31260 61152 31305 61180
rect 31260 61140 31266 61152
rect 31665 61149 31677 61183
rect 31711 61180 31723 61183
rect 31754 61180 31760 61192
rect 31711 61152 31760 61180
rect 31711 61149 31723 61152
rect 31665 61143 31723 61149
rect 31754 61140 31760 61152
rect 31812 61180 31818 61192
rect 32398 61180 32404 61192
rect 31812 61152 32404 61180
rect 31812 61140 31818 61152
rect 32398 61140 32404 61152
rect 32456 61140 32462 61192
rect 34698 61140 34704 61192
rect 34756 61180 34762 61192
rect 34977 61183 35035 61189
rect 34977 61180 34989 61183
rect 34756 61152 34989 61180
rect 34756 61140 34762 61152
rect 34977 61149 34989 61152
rect 35023 61149 35035 61183
rect 34977 61143 35035 61149
rect 35066 61140 35072 61192
rect 35124 61180 35130 61192
rect 35342 61180 35348 61192
rect 35124 61152 35348 61180
rect 35124 61140 35130 61152
rect 35342 61140 35348 61152
rect 35400 61140 35406 61192
rect 35986 61180 35992 61192
rect 35947 61152 35992 61180
rect 35986 61140 35992 61152
rect 36044 61140 36050 61192
rect 36096 61189 36124 61276
rect 36081 61183 36139 61189
rect 36081 61149 36093 61183
rect 36127 61149 36139 61183
rect 36081 61143 36139 61149
rect 36170 61140 36176 61192
rect 36228 61180 36234 61192
rect 36354 61180 36360 61192
rect 36228 61152 36273 61180
rect 36315 61152 36360 61180
rect 36228 61140 36234 61152
rect 36354 61140 36360 61152
rect 36412 61140 36418 61192
rect 36832 61189 36860 61356
rect 67634 61344 67640 61356
rect 67692 61344 67698 61396
rect 36817 61183 36875 61189
rect 36817 61149 36829 61183
rect 36863 61180 36875 61183
rect 37366 61180 37372 61192
rect 36863 61152 37372 61180
rect 36863 61149 36875 61152
rect 36817 61143 36875 61149
rect 37366 61140 37372 61152
rect 37424 61180 37430 61192
rect 38102 61180 38108 61192
rect 37424 61152 38108 61180
rect 37424 61140 37430 61152
rect 38102 61140 38108 61152
rect 38160 61180 38166 61192
rect 38933 61183 38991 61189
rect 38933 61180 38945 61183
rect 38160 61152 38945 61180
rect 38160 61140 38166 61152
rect 38933 61149 38945 61152
rect 38979 61180 38991 61183
rect 39853 61183 39911 61189
rect 39853 61180 39865 61183
rect 38979 61152 39865 61180
rect 38979 61149 38991 61152
rect 38933 61143 38991 61149
rect 39853 61149 39865 61152
rect 39899 61180 39911 61183
rect 39942 61180 39948 61192
rect 39899 61152 39948 61180
rect 39899 61149 39911 61152
rect 39853 61143 39911 61149
rect 39942 61140 39948 61152
rect 40000 61140 40006 61192
rect 67542 61180 67548 61192
rect 67503 61152 67548 61180
rect 67542 61140 67548 61152
rect 67600 61140 67606 61192
rect 28368 61112 28396 61140
rect 27540 61084 28396 61112
rect 30561 61115 30619 61121
rect 30561 61081 30573 61115
rect 30607 61112 30619 61115
rect 31910 61115 31968 61121
rect 31910 61112 31922 61115
rect 30607 61084 31922 61112
rect 30607 61081 30619 61084
rect 30561 61075 30619 61081
rect 31910 61081 31922 61084
rect 31956 61081 31968 61115
rect 31910 61075 31968 61081
rect 34793 61115 34851 61121
rect 34793 61081 34805 61115
rect 34839 61112 34851 61115
rect 35526 61112 35532 61124
rect 34839 61084 35532 61112
rect 34839 61081 34851 61084
rect 34793 61075 34851 61081
rect 35526 61072 35532 61084
rect 35584 61072 35590 61124
rect 37062 61115 37120 61121
rect 37062 61112 37074 61115
rect 36280 61084 37074 61112
rect 20806 61044 20812 61056
rect 20272 61016 20812 61044
rect 20806 61004 20812 61016
rect 20864 61044 20870 61056
rect 22557 61047 22615 61053
rect 22557 61044 22569 61047
rect 20864 61016 22569 61044
rect 20864 61004 20870 61016
rect 22557 61013 22569 61016
rect 22603 61013 22615 61047
rect 22557 61007 22615 61013
rect 35713 61047 35771 61053
rect 35713 61013 35725 61047
rect 35759 61044 35771 61047
rect 36280 61044 36308 61084
rect 37062 61081 37074 61084
rect 37108 61081 37120 61115
rect 38746 61112 38752 61124
rect 38707 61084 38752 61112
rect 37062 61075 37120 61081
rect 38746 61072 38752 61084
rect 38804 61072 38810 61124
rect 40126 61121 40132 61124
rect 40120 61075 40132 61121
rect 40184 61112 40190 61124
rect 40184 61084 40220 61112
rect 40126 61072 40132 61075
rect 40184 61072 40190 61084
rect 35759 61016 36308 61044
rect 35759 61013 35771 61016
rect 35713 61007 35771 61013
rect 36538 61004 36544 61056
rect 36596 61044 36602 61056
rect 38197 61047 38255 61053
rect 38197 61044 38209 61047
rect 36596 61016 38209 61044
rect 36596 61004 36602 61016
rect 38197 61013 38209 61016
rect 38243 61013 38255 61047
rect 41230 61044 41236 61056
rect 41191 61016 41236 61044
rect 38197 61007 38255 61013
rect 41230 61004 41236 61016
rect 41288 61004 41294 61056
rect 1104 60954 68816 60976
rect 1104 60902 19574 60954
rect 19626 60902 19638 60954
rect 19690 60902 19702 60954
rect 19754 60902 19766 60954
rect 19818 60902 19830 60954
rect 19882 60902 50294 60954
rect 50346 60902 50358 60954
rect 50410 60902 50422 60954
rect 50474 60902 50486 60954
rect 50538 60902 50550 60954
rect 50602 60902 68816 60954
rect 1104 60880 68816 60902
rect 19334 60800 19340 60852
rect 19392 60840 19398 60852
rect 19521 60843 19579 60849
rect 19521 60840 19533 60843
rect 19392 60812 19533 60840
rect 19392 60800 19398 60812
rect 19521 60809 19533 60812
rect 19567 60809 19579 60843
rect 19521 60803 19579 60809
rect 26234 60800 26240 60852
rect 26292 60840 26298 60852
rect 30282 60840 30288 60852
rect 26292 60812 26337 60840
rect 30243 60812 30288 60840
rect 26292 60800 26298 60812
rect 30282 60800 30288 60812
rect 30340 60800 30346 60852
rect 36354 60800 36360 60852
rect 36412 60840 36418 60852
rect 36633 60843 36691 60849
rect 36633 60840 36645 60843
rect 36412 60812 36645 60840
rect 36412 60800 36418 60812
rect 36633 60809 36645 60812
rect 36679 60809 36691 60843
rect 36633 60803 36691 60809
rect 40037 60843 40095 60849
rect 40037 60809 40049 60843
rect 40083 60840 40095 60843
rect 40126 60840 40132 60852
rect 40083 60812 40132 60840
rect 40083 60809 40095 60812
rect 40037 60803 40095 60809
rect 40126 60800 40132 60812
rect 40184 60800 40190 60852
rect 1854 60772 1860 60784
rect 1815 60744 1860 60772
rect 1854 60732 1860 60744
rect 1912 60732 1918 60784
rect 31478 60772 31484 60784
rect 30668 60744 31484 60772
rect 16117 60707 16175 60713
rect 16117 60673 16129 60707
rect 16163 60704 16175 60707
rect 17034 60704 17040 60716
rect 16163 60676 17040 60704
rect 16163 60673 16175 60676
rect 16117 60667 16175 60673
rect 17034 60664 17040 60676
rect 17092 60664 17098 60716
rect 17494 60664 17500 60716
rect 17552 60704 17558 60716
rect 17661 60707 17719 60713
rect 17661 60704 17673 60707
rect 17552 60676 17673 60704
rect 17552 60664 17558 60676
rect 17661 60673 17673 60676
rect 17707 60673 17719 60707
rect 17661 60667 17719 60673
rect 19705 60707 19763 60713
rect 19705 60673 19717 60707
rect 19751 60704 19763 60707
rect 19978 60704 19984 60716
rect 19751 60676 19984 60704
rect 19751 60673 19763 60676
rect 19705 60667 19763 60673
rect 19978 60664 19984 60676
rect 20036 60664 20042 60716
rect 22373 60707 22431 60713
rect 22373 60704 22385 60707
rect 20088 60676 22385 60704
rect 17402 60636 17408 60648
rect 17363 60608 17408 60636
rect 17402 60596 17408 60608
rect 17460 60596 17466 60648
rect 20088 60568 20116 60676
rect 22373 60673 22385 60676
rect 22419 60673 22431 60707
rect 22373 60667 22431 60673
rect 23477 60707 23535 60713
rect 23477 60673 23489 60707
rect 23523 60673 23535 60707
rect 23477 60667 23535 60673
rect 25133 60707 25191 60713
rect 25133 60673 25145 60707
rect 25179 60704 25191 60707
rect 25498 60704 25504 60716
rect 25179 60676 25504 60704
rect 25179 60673 25191 60676
rect 25133 60667 25191 60673
rect 22002 60596 22008 60648
rect 22060 60636 22066 60648
rect 22189 60639 22247 60645
rect 22189 60636 22201 60639
rect 22060 60608 22201 60636
rect 22060 60596 22066 60608
rect 22189 60605 22201 60608
rect 22235 60605 22247 60639
rect 23492 60636 23520 60667
rect 25498 60664 25504 60676
rect 25556 60664 25562 60716
rect 26421 60707 26479 60713
rect 26421 60673 26433 60707
rect 26467 60704 26479 60707
rect 27433 60707 27491 60713
rect 26467 60676 27384 60704
rect 26467 60673 26479 60676
rect 26421 60667 26479 60673
rect 26326 60636 26332 60648
rect 23492 60608 26332 60636
rect 22189 60599 22247 60605
rect 26326 60596 26332 60608
rect 26384 60596 26390 60648
rect 27249 60639 27307 60645
rect 27249 60605 27261 60639
rect 27295 60605 27307 60639
rect 27356 60636 27384 60676
rect 27433 60673 27445 60707
rect 27479 60704 27491 60707
rect 27706 60704 27712 60716
rect 27479 60676 27712 60704
rect 27479 60673 27491 60676
rect 27433 60667 27491 60673
rect 27706 60664 27712 60676
rect 27764 60664 27770 60716
rect 30374 60664 30380 60716
rect 30432 60704 30438 60716
rect 30668 60713 30696 60744
rect 31478 60732 31484 60744
rect 31536 60732 31542 60784
rect 30561 60707 30619 60713
rect 30561 60704 30573 60707
rect 30432 60676 30573 60704
rect 30432 60664 30438 60676
rect 30561 60673 30573 60676
rect 30607 60673 30619 60707
rect 30561 60667 30619 60673
rect 30653 60707 30711 60713
rect 30653 60673 30665 60707
rect 30699 60704 30711 60707
rect 30766 60707 30824 60713
rect 30699 60676 30733 60704
rect 30699 60673 30711 60676
rect 30653 60667 30711 60673
rect 30766 60673 30778 60707
rect 30812 60704 30824 60707
rect 30929 60707 30987 60713
rect 30812 60676 30880 60704
rect 30812 60673 30824 60676
rect 30766 60667 30824 60673
rect 27617 60639 27675 60645
rect 27617 60636 27629 60639
rect 27356 60608 27629 60636
rect 27249 60599 27307 60605
rect 27617 60605 27629 60608
rect 27663 60605 27675 60639
rect 27617 60599 27675 60605
rect 18340 60540 20116 60568
rect 2130 60500 2136 60512
rect 2091 60472 2136 60500
rect 2130 60460 2136 60472
rect 2188 60460 2194 60512
rect 15838 60460 15844 60512
rect 15896 60500 15902 60512
rect 15933 60503 15991 60509
rect 15933 60500 15945 60503
rect 15896 60472 15945 60500
rect 15896 60460 15902 60472
rect 15933 60469 15945 60472
rect 15979 60469 15991 60503
rect 15933 60463 15991 60469
rect 16022 60460 16028 60512
rect 16080 60500 16086 60512
rect 18340 60500 18368 60540
rect 23658 60528 23664 60580
rect 23716 60568 23722 60580
rect 27264 60568 27292 60599
rect 30466 60596 30472 60648
rect 30524 60636 30530 60648
rect 30852 60636 30880 60676
rect 30929 60673 30941 60707
rect 30975 60704 30987 60707
rect 31202 60704 31208 60716
rect 30975 60676 31208 60704
rect 30975 60673 30987 60676
rect 30929 60667 30987 60673
rect 30524 60608 30880 60636
rect 30524 60596 30530 60608
rect 28074 60568 28080 60580
rect 23716 60540 25084 60568
rect 27264 60540 28080 60568
rect 23716 60528 23722 60540
rect 18782 60500 18788 60512
rect 16080 60472 18368 60500
rect 18695 60472 18788 60500
rect 16080 60460 16086 60472
rect 18782 60460 18788 60472
rect 18840 60500 18846 60512
rect 21542 60500 21548 60512
rect 18840 60472 21548 60500
rect 18840 60460 18846 60472
rect 21542 60460 21548 60472
rect 21600 60460 21606 60512
rect 22370 60460 22376 60512
rect 22428 60500 22434 60512
rect 22557 60503 22615 60509
rect 22557 60500 22569 60503
rect 22428 60472 22569 60500
rect 22428 60460 22434 60472
rect 22557 60469 22569 60472
rect 22603 60469 22615 60503
rect 22557 60463 22615 60469
rect 22830 60460 22836 60512
rect 22888 60500 22894 60512
rect 23569 60503 23627 60509
rect 23569 60500 23581 60503
rect 22888 60472 23581 60500
rect 22888 60460 22894 60472
rect 23569 60469 23581 60472
rect 23615 60469 23627 60503
rect 24946 60500 24952 60512
rect 24907 60472 24952 60500
rect 23569 60463 23627 60469
rect 24946 60460 24952 60472
rect 25004 60460 25010 60512
rect 25056 60500 25084 60540
rect 28074 60528 28080 60540
rect 28132 60528 28138 60580
rect 30944 60500 30972 60667
rect 31202 60664 31208 60676
rect 31260 60664 31266 60716
rect 33686 60704 33692 60716
rect 33647 60676 33692 60704
rect 33686 60664 33692 60676
rect 33744 60664 33750 60716
rect 35897 60707 35955 60713
rect 35897 60673 35909 60707
rect 35943 60704 35955 60707
rect 36078 60704 36084 60716
rect 35943 60676 36084 60704
rect 35943 60673 35955 60676
rect 35897 60667 35955 60673
rect 36078 60664 36084 60676
rect 36136 60704 36142 60716
rect 36538 60704 36544 60716
rect 36136 60676 36544 60704
rect 36136 60664 36142 60676
rect 36538 60664 36544 60676
rect 36596 60664 36602 60716
rect 36725 60707 36783 60713
rect 36725 60673 36737 60707
rect 36771 60673 36783 60707
rect 38102 60704 38108 60716
rect 38063 60676 38108 60704
rect 36725 60667 36783 60673
rect 35713 60639 35771 60645
rect 35713 60605 35725 60639
rect 35759 60636 35771 60639
rect 35986 60636 35992 60648
rect 35759 60608 35992 60636
rect 35759 60605 35771 60608
rect 35713 60599 35771 60605
rect 35986 60596 35992 60608
rect 36044 60636 36050 60648
rect 36740 60636 36768 60667
rect 38102 60664 38108 60676
rect 38160 60664 38166 60716
rect 38372 60707 38430 60713
rect 38372 60673 38384 60707
rect 38418 60704 38430 60707
rect 38654 60704 38660 60716
rect 38418 60676 38660 60704
rect 38418 60673 38430 60676
rect 38372 60667 38430 60673
rect 38654 60664 38660 60676
rect 38712 60664 38718 60716
rect 39850 60664 39856 60716
rect 39908 60704 39914 60716
rect 39945 60707 40003 60713
rect 39945 60704 39957 60707
rect 39908 60676 39957 60704
rect 39908 60664 39914 60676
rect 39945 60673 39957 60676
rect 39991 60673 40003 60707
rect 40126 60704 40132 60716
rect 40087 60676 40132 60704
rect 39945 60667 40003 60673
rect 40126 60664 40132 60676
rect 40184 60664 40190 60716
rect 36044 60608 36768 60636
rect 65797 60639 65855 60645
rect 36044 60596 36050 60608
rect 65797 60605 65809 60639
rect 65843 60605 65855 60639
rect 65797 60599 65855 60605
rect 65981 60639 66039 60645
rect 65981 60605 65993 60639
rect 66027 60636 66039 60639
rect 67358 60636 67364 60648
rect 66027 60608 67364 60636
rect 66027 60605 66039 60608
rect 65981 60599 66039 60605
rect 35066 60528 35072 60580
rect 35124 60568 35130 60580
rect 36081 60571 36139 60577
rect 36081 60568 36093 60571
rect 35124 60540 36093 60568
rect 35124 60528 35130 60540
rect 36081 60537 36093 60540
rect 36127 60537 36139 60571
rect 65812 60568 65840 60599
rect 67358 60596 67364 60608
rect 67416 60596 67422 60648
rect 67542 60636 67548 60648
rect 67503 60608 67548 60636
rect 67542 60596 67548 60608
rect 67600 60596 67606 60648
rect 68094 60568 68100 60580
rect 65812 60540 68100 60568
rect 36081 60531 36139 60537
rect 68094 60528 68100 60540
rect 68152 60528 68158 60580
rect 25056 60472 30972 60500
rect 33781 60503 33839 60509
rect 33781 60469 33793 60503
rect 33827 60500 33839 60503
rect 33962 60500 33968 60512
rect 33827 60472 33968 60500
rect 33827 60469 33839 60472
rect 33781 60463 33839 60469
rect 33962 60460 33968 60472
rect 34020 60460 34026 60512
rect 39206 60460 39212 60512
rect 39264 60500 39270 60512
rect 39485 60503 39543 60509
rect 39485 60500 39497 60503
rect 39264 60472 39497 60500
rect 39264 60460 39270 60472
rect 39485 60469 39497 60472
rect 39531 60469 39543 60503
rect 39485 60463 39543 60469
rect 1104 60410 68816 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 65654 60410
rect 65706 60358 65718 60410
rect 65770 60358 65782 60410
rect 65834 60358 65846 60410
rect 65898 60358 65910 60410
rect 65962 60358 68816 60410
rect 1104 60336 68816 60358
rect 19978 60256 19984 60308
rect 20036 60296 20042 60308
rect 20036 60268 25728 60296
rect 20036 60256 20042 60268
rect 19242 60188 19248 60240
rect 19300 60228 19306 60240
rect 21453 60231 21511 60237
rect 21453 60228 21465 60231
rect 19300 60200 21465 60228
rect 19300 60188 19306 60200
rect 21453 60197 21465 60200
rect 21499 60197 21511 60231
rect 21453 60191 21511 60197
rect 17405 60163 17463 60169
rect 17405 60129 17417 60163
rect 17451 60160 17463 60163
rect 18782 60160 18788 60172
rect 17451 60132 18788 60160
rect 17451 60129 17463 60132
rect 17405 60123 17463 60129
rect 18782 60120 18788 60132
rect 18840 60120 18846 60172
rect 20806 60160 20812 60172
rect 20767 60132 20812 60160
rect 20806 60120 20812 60132
rect 20864 60120 20870 60172
rect 21542 60120 21548 60172
rect 21600 60160 21606 60172
rect 21846 60163 21904 60169
rect 21846 60160 21858 60163
rect 21600 60132 21858 60160
rect 21600 60120 21606 60132
rect 21846 60129 21858 60132
rect 21892 60129 21904 60163
rect 21846 60123 21904 60129
rect 22005 60163 22063 60169
rect 22005 60129 22017 60163
rect 22051 60160 22063 60163
rect 22388 60160 22416 60268
rect 25700 60228 25728 60268
rect 25774 60256 25780 60308
rect 25832 60296 25838 60308
rect 28258 60296 28264 60308
rect 25832 60268 28264 60296
rect 25832 60256 25838 60268
rect 28258 60256 28264 60268
rect 28316 60256 28322 60308
rect 30377 60299 30435 60305
rect 30377 60265 30389 60299
rect 30423 60296 30435 60299
rect 30466 60296 30472 60308
rect 30423 60268 30472 60296
rect 30423 60265 30435 60268
rect 30377 60259 30435 60265
rect 30466 60256 30472 60268
rect 30524 60256 30530 60308
rect 31018 60256 31024 60308
rect 31076 60296 31082 60308
rect 31297 60299 31355 60305
rect 31297 60296 31309 60299
rect 31076 60268 31309 60296
rect 31076 60256 31082 60268
rect 31297 60265 31309 60268
rect 31343 60265 31355 60299
rect 31297 60259 31355 60265
rect 38654 60256 38660 60308
rect 38712 60296 38718 60308
rect 38749 60299 38807 60305
rect 38749 60296 38761 60299
rect 38712 60268 38761 60296
rect 38712 60256 38718 60268
rect 38749 60265 38761 60268
rect 38795 60265 38807 60299
rect 38749 60259 38807 60265
rect 39853 60299 39911 60305
rect 39853 60265 39865 60299
rect 39899 60296 39911 60299
rect 40126 60296 40132 60308
rect 39899 60268 40132 60296
rect 39899 60265 39911 60268
rect 39853 60259 39911 60265
rect 40126 60256 40132 60268
rect 40184 60256 40190 60308
rect 67358 60296 67364 60308
rect 67319 60268 67364 60296
rect 67358 60256 67364 60268
rect 67416 60256 67422 60308
rect 68094 60296 68100 60308
rect 68055 60268 68100 60296
rect 68094 60256 68100 60268
rect 68152 60256 68158 60308
rect 27614 60228 27620 60240
rect 25700 60200 27620 60228
rect 27614 60188 27620 60200
rect 27672 60188 27678 60240
rect 22051 60132 22416 60160
rect 27157 60163 27215 60169
rect 22051 60129 22063 60132
rect 22005 60123 22063 60129
rect 27157 60129 27169 60163
rect 27203 60160 27215 60163
rect 27430 60160 27436 60172
rect 27203 60132 27436 60160
rect 27203 60129 27215 60132
rect 27157 60123 27215 60129
rect 27430 60120 27436 60132
rect 27488 60120 27494 60172
rect 27798 60160 27804 60172
rect 27759 60132 27804 60160
rect 27798 60120 27804 60132
rect 27856 60120 27862 60172
rect 28258 60169 28264 60172
rect 28215 60163 28264 60169
rect 28215 60129 28227 60163
rect 28261 60129 28264 60163
rect 28215 60123 28264 60129
rect 28258 60120 28264 60123
rect 28316 60120 28322 60172
rect 28534 60160 28540 60172
rect 28368 60132 28540 60160
rect 1670 60052 1676 60104
rect 1728 60092 1734 60104
rect 1857 60095 1915 60101
rect 1857 60092 1869 60095
rect 1728 60064 1869 60092
rect 1728 60052 1734 60064
rect 1857 60061 1869 60064
rect 1903 60061 1915 60095
rect 15562 60092 15568 60104
rect 15523 60064 15568 60092
rect 1857 60055 1915 60061
rect 15562 60052 15568 60064
rect 15620 60052 15626 60104
rect 15838 60101 15844 60104
rect 15832 60092 15844 60101
rect 15799 60064 15844 60092
rect 15832 60055 15844 60064
rect 15838 60052 15844 60055
rect 15896 60052 15902 60104
rect 16574 60052 16580 60104
rect 16632 60092 16638 60104
rect 17589 60095 17647 60101
rect 17589 60092 17601 60095
rect 16632 60064 17601 60092
rect 16632 60052 16638 60064
rect 17589 60061 17601 60064
rect 17635 60061 17647 60095
rect 20990 60092 20996 60104
rect 20951 60064 20996 60092
rect 17589 60055 17647 60061
rect 20990 60052 20996 60064
rect 21048 60052 21054 60104
rect 21726 60052 21732 60104
rect 21784 60092 21790 60104
rect 23750 60092 23756 60104
rect 21784 60064 21829 60092
rect 23711 60064 23756 60092
rect 21784 60052 21790 60064
rect 23750 60052 23756 60064
rect 23808 60052 23814 60104
rect 23845 60095 23903 60101
rect 23845 60061 23857 60095
rect 23891 60092 23903 60095
rect 24397 60095 24455 60101
rect 24397 60092 24409 60095
rect 23891 60064 24409 60092
rect 23891 60061 23903 60064
rect 23845 60055 23903 60061
rect 24397 60061 24409 60064
rect 24443 60061 24455 60095
rect 24397 60055 24455 60061
rect 24664 60095 24722 60101
rect 24664 60061 24676 60095
rect 24710 60092 24722 60095
rect 24946 60092 24952 60104
rect 24710 60064 24952 60092
rect 24710 60061 24722 60064
rect 24664 60055 24722 60061
rect 24946 60052 24952 60064
rect 25004 60052 25010 60104
rect 26326 60092 26332 60104
rect 26287 60064 26332 60092
rect 26326 60052 26332 60064
rect 26384 60052 26390 60104
rect 27341 60095 27399 60101
rect 27341 60061 27353 60095
rect 27387 60061 27399 60095
rect 27341 60055 27399 60061
rect 23768 60024 23796 60052
rect 22572 59996 23796 60024
rect 16942 59956 16948 59968
rect 16903 59928 16948 59956
rect 16942 59916 16948 59928
rect 17000 59916 17006 59968
rect 17586 59916 17592 59968
rect 17644 59956 17650 59968
rect 17773 59959 17831 59965
rect 17773 59956 17785 59959
rect 17644 59928 17785 59956
rect 17644 59916 17650 59928
rect 17773 59925 17785 59928
rect 17819 59925 17831 59959
rect 17773 59919 17831 59925
rect 17862 59916 17868 59968
rect 17920 59956 17926 59968
rect 22572 59956 22600 59996
rect 17920 59928 22600 59956
rect 22649 59959 22707 59965
rect 17920 59916 17926 59928
rect 22649 59925 22661 59959
rect 22695 59956 22707 59959
rect 26326 59956 26332 59968
rect 22695 59928 26332 59956
rect 22695 59925 22707 59928
rect 22649 59919 22707 59925
rect 26326 59916 26332 59928
rect 26384 59916 26390 59968
rect 26421 59959 26479 59965
rect 26421 59925 26433 59959
rect 26467 59956 26479 59959
rect 26970 59956 26976 59968
rect 26467 59928 26976 59956
rect 26467 59925 26479 59928
rect 26421 59919 26479 59925
rect 26970 59916 26976 59928
rect 27028 59916 27034 59968
rect 27356 59956 27384 60055
rect 28074 60052 28080 60104
rect 28132 60092 28138 60104
rect 28368 60101 28396 60132
rect 28534 60120 28540 60132
rect 28592 60120 28598 60172
rect 30576 60132 31524 60160
rect 28353 60095 28411 60101
rect 28132 60064 28177 60092
rect 28132 60052 28138 60064
rect 28353 60061 28365 60095
rect 28399 60061 28411 60095
rect 28353 60055 28411 60061
rect 29733 60095 29791 60101
rect 29733 60061 29745 60095
rect 29779 60092 29791 60095
rect 29914 60092 29920 60104
rect 29779 60064 29920 60092
rect 29779 60061 29791 60064
rect 29733 60055 29791 60061
rect 29914 60052 29920 60064
rect 29972 60052 29978 60104
rect 30576 60101 30604 60132
rect 31496 60101 31524 60132
rect 38838 60120 38844 60172
rect 38896 60160 38902 60172
rect 39117 60163 39175 60169
rect 39117 60160 39129 60163
rect 38896 60132 39129 60160
rect 38896 60120 38902 60132
rect 39117 60129 39129 60132
rect 39163 60129 39175 60163
rect 39117 60123 39175 60129
rect 39942 60120 39948 60172
rect 40000 60160 40006 60172
rect 42889 60163 42947 60169
rect 42889 60160 42901 60163
rect 40000 60132 42901 60160
rect 40000 60120 40006 60132
rect 42889 60129 42901 60132
rect 42935 60129 42947 60163
rect 42889 60123 42947 60129
rect 30561 60095 30619 60101
rect 30561 60061 30573 60095
rect 30607 60061 30619 60095
rect 30561 60055 30619 60061
rect 30837 60095 30895 60101
rect 30837 60061 30849 60095
rect 30883 60061 30895 60095
rect 30837 60055 30895 60061
rect 31481 60095 31539 60101
rect 31481 60061 31493 60095
rect 31527 60092 31539 60095
rect 31662 60092 31668 60104
rect 31527 60064 31668 60092
rect 31527 60061 31539 60064
rect 31481 60055 31539 60061
rect 28997 60027 29055 60033
rect 28997 59993 29009 60027
rect 29043 60024 29055 60027
rect 30852 60024 30880 60055
rect 31662 60052 31668 60064
rect 31720 60052 31726 60104
rect 31754 60052 31760 60104
rect 31812 60092 31818 60104
rect 31812 60064 31857 60092
rect 31812 60052 31818 60064
rect 32398 60052 32404 60104
rect 32456 60092 32462 60104
rect 32677 60095 32735 60101
rect 32677 60092 32689 60095
rect 32456 60064 32689 60092
rect 32456 60052 32462 60064
rect 32677 60061 32689 60064
rect 32723 60092 32735 60095
rect 35529 60095 35587 60101
rect 32723 60064 33088 60092
rect 32723 60061 32735 60064
rect 32677 60055 32735 60061
rect 33060 60036 33088 60064
rect 35529 60061 35541 60095
rect 35575 60092 35587 60095
rect 36538 60092 36544 60104
rect 35575 60064 36544 60092
rect 35575 60061 35587 60064
rect 35529 60055 35587 60061
rect 36538 60052 36544 60064
rect 36596 60052 36602 60104
rect 38930 60092 38936 60104
rect 38891 60064 38936 60092
rect 38930 60052 38936 60064
rect 38988 60052 38994 60104
rect 39209 60095 39267 60101
rect 39209 60061 39221 60095
rect 39255 60092 39267 60095
rect 39666 60092 39672 60104
rect 39255 60064 39672 60092
rect 39255 60061 39267 60064
rect 39209 60055 39267 60061
rect 39666 60052 39672 60064
rect 39724 60092 39730 60104
rect 40037 60095 40095 60101
rect 40037 60092 40049 60095
rect 39724 60064 40049 60092
rect 39724 60052 39730 60064
rect 40037 60061 40049 60064
rect 40083 60061 40095 60095
rect 40037 60055 40095 60061
rect 40126 60052 40132 60104
rect 40184 60092 40190 60104
rect 40184 60064 40229 60092
rect 40184 60052 40190 60064
rect 42702 60052 42708 60104
rect 42760 60092 42766 60104
rect 67269 60095 67327 60101
rect 67269 60092 67281 60095
rect 42760 60064 67281 60092
rect 42760 60052 42766 60064
rect 67269 60061 67281 60064
rect 67315 60061 67327 60095
rect 67269 60055 67327 60061
rect 29043 59996 30880 60024
rect 29043 59993 29055 59996
rect 28997 59987 29055 59993
rect 32214 59984 32220 60036
rect 32272 60024 32278 60036
rect 32922 60027 32980 60033
rect 32922 60024 32934 60027
rect 32272 59996 32934 60024
rect 32272 59984 32278 59996
rect 32922 59993 32934 59996
rect 32968 59993 32980 60027
rect 32922 59987 32980 59993
rect 33042 59984 33048 60036
rect 33100 59984 33106 60036
rect 39853 60027 39911 60033
rect 39853 59993 39865 60027
rect 39899 60024 39911 60027
rect 40218 60024 40224 60036
rect 39899 59996 40224 60024
rect 39899 59993 39911 59996
rect 39853 59987 39911 59993
rect 40218 59984 40224 59996
rect 40276 60024 40282 60036
rect 41230 60024 41236 60036
rect 40276 59996 41236 60024
rect 40276 59984 40282 59996
rect 41230 59984 41236 59996
rect 41288 59984 41294 60036
rect 43156 60027 43214 60033
rect 43156 59993 43168 60027
rect 43202 60024 43214 60027
rect 44082 60024 44088 60036
rect 43202 59996 44088 60024
rect 43202 59993 43214 59996
rect 43156 59987 43214 59993
rect 44082 59984 44088 59996
rect 44140 59984 44146 60036
rect 29270 59956 29276 59968
rect 27356 59928 29276 59956
rect 29270 59916 29276 59928
rect 29328 59916 29334 59968
rect 29549 59959 29607 59965
rect 29549 59925 29561 59959
rect 29595 59956 29607 59959
rect 29638 59956 29644 59968
rect 29595 59928 29644 59956
rect 29595 59925 29607 59928
rect 29549 59919 29607 59925
rect 29638 59916 29644 59928
rect 29696 59916 29702 59968
rect 30745 59959 30803 59965
rect 30745 59925 30757 59959
rect 30791 59956 30803 59959
rect 31665 59959 31723 59965
rect 31665 59956 31677 59959
rect 30791 59928 31677 59956
rect 30791 59925 30803 59928
rect 30745 59919 30803 59925
rect 31665 59925 31677 59928
rect 31711 59956 31723 59959
rect 31846 59956 31852 59968
rect 31711 59928 31852 59956
rect 31711 59925 31723 59928
rect 31665 59919 31723 59925
rect 31846 59916 31852 59928
rect 31904 59916 31910 59968
rect 33778 59916 33784 59968
rect 33836 59956 33842 59968
rect 34057 59959 34115 59965
rect 34057 59956 34069 59959
rect 33836 59928 34069 59956
rect 33836 59916 33842 59928
rect 34057 59925 34069 59928
rect 34103 59925 34115 59959
rect 35342 59956 35348 59968
rect 35303 59928 35348 59956
rect 34057 59919 34115 59925
rect 35342 59916 35348 59928
rect 35400 59916 35406 59968
rect 42978 59916 42984 59968
rect 43036 59956 43042 59968
rect 44269 59959 44327 59965
rect 44269 59956 44281 59959
rect 43036 59928 44281 59956
rect 43036 59916 43042 59928
rect 44269 59925 44281 59928
rect 44315 59925 44327 59959
rect 44269 59919 44327 59925
rect 1104 59866 68816 59888
rect 1104 59814 19574 59866
rect 19626 59814 19638 59866
rect 19690 59814 19702 59866
rect 19754 59814 19766 59866
rect 19818 59814 19830 59866
rect 19882 59814 50294 59866
rect 50346 59814 50358 59866
rect 50410 59814 50422 59866
rect 50474 59814 50486 59866
rect 50538 59814 50550 59866
rect 50602 59814 68816 59866
rect 1104 59792 68816 59814
rect 15562 59712 15568 59764
rect 15620 59752 15626 59764
rect 15841 59755 15899 59761
rect 15841 59752 15853 59755
rect 15620 59724 15853 59752
rect 15620 59712 15626 59724
rect 15841 59721 15853 59724
rect 15887 59721 15899 59755
rect 17034 59752 17040 59764
rect 16995 59724 17040 59752
rect 15841 59715 15899 59721
rect 17034 59712 17040 59724
rect 17092 59712 17098 59764
rect 17402 59712 17408 59764
rect 17460 59752 17466 59764
rect 17681 59755 17739 59761
rect 17681 59752 17693 59755
rect 17460 59724 17693 59752
rect 17460 59712 17466 59724
rect 17681 59721 17693 59724
rect 17727 59721 17739 59755
rect 19426 59752 19432 59764
rect 17681 59715 17739 59721
rect 18708 59724 19432 59752
rect 15856 59656 17724 59684
rect 15856 59628 15884 59656
rect 1670 59616 1676 59628
rect 1631 59588 1676 59616
rect 1670 59576 1676 59588
rect 1728 59576 1734 59628
rect 14642 59616 14648 59628
rect 14603 59588 14648 59616
rect 14642 59576 14648 59588
rect 14700 59576 14706 59628
rect 15838 59616 15844 59628
rect 15751 59588 15844 59616
rect 15838 59576 15844 59588
rect 15896 59576 15902 59628
rect 16574 59576 16580 59628
rect 16632 59616 16638 59628
rect 17696 59625 17724 59656
rect 16853 59619 16911 59625
rect 16853 59616 16865 59619
rect 16632 59588 16865 59616
rect 16632 59576 16638 59588
rect 16853 59585 16865 59588
rect 16899 59585 16911 59619
rect 16853 59579 16911 59585
rect 17681 59619 17739 59625
rect 17681 59585 17693 59619
rect 17727 59616 17739 59619
rect 17862 59616 17868 59628
rect 17727 59588 17868 59616
rect 17727 59585 17739 59588
rect 17681 59579 17739 59585
rect 17862 59576 17868 59588
rect 17920 59576 17926 59628
rect 18601 59619 18659 59625
rect 18601 59585 18613 59619
rect 18647 59616 18659 59619
rect 18708 59616 18736 59724
rect 19426 59712 19432 59724
rect 19484 59712 19490 59764
rect 22189 59755 22247 59761
rect 22189 59721 22201 59755
rect 22235 59721 22247 59755
rect 25498 59752 25504 59764
rect 25459 59724 25504 59752
rect 22189 59715 22247 59721
rect 22204 59684 22232 59715
rect 25498 59712 25504 59724
rect 25556 59712 25562 59764
rect 26326 59712 26332 59764
rect 26384 59752 26390 59764
rect 26384 59724 27384 59752
rect 26384 59712 26390 59724
rect 23078 59687 23136 59693
rect 23078 59684 23090 59687
rect 22204 59656 23090 59684
rect 23078 59653 23090 59656
rect 23124 59653 23136 59687
rect 25774 59684 25780 59696
rect 23078 59647 23136 59653
rect 25240 59656 25780 59684
rect 18647 59588 18736 59616
rect 18647 59585 18659 59588
rect 18601 59579 18659 59585
rect 18782 59576 18788 59628
rect 18840 59616 18846 59628
rect 18840 59588 18885 59616
rect 18840 59576 18846 59588
rect 19518 59576 19524 59628
rect 19576 59616 19582 59628
rect 22370 59616 22376 59628
rect 19576 59588 19621 59616
rect 22331 59588 22376 59616
rect 19576 59576 19582 59588
rect 22370 59576 22376 59588
rect 22428 59576 22434 59628
rect 22830 59616 22836 59628
rect 22791 59588 22836 59616
rect 22830 59576 22836 59588
rect 22888 59576 22894 59628
rect 25240 59625 25268 59656
rect 25774 59644 25780 59656
rect 25832 59644 25838 59696
rect 26234 59644 26240 59696
rect 26292 59684 26298 59696
rect 27218 59687 27276 59693
rect 27218 59684 27230 59687
rect 26292 59656 27230 59684
rect 26292 59644 26298 59656
rect 27218 59653 27230 59656
rect 27264 59653 27276 59687
rect 27356 59684 27384 59724
rect 28074 59712 28080 59764
rect 28132 59752 28138 59764
rect 28353 59755 28411 59761
rect 28353 59752 28365 59755
rect 28132 59724 28365 59752
rect 28132 59712 28138 59724
rect 28353 59721 28365 59724
rect 28399 59721 28411 59755
rect 32214 59752 32220 59764
rect 32175 59724 32220 59752
rect 28353 59715 28411 59721
rect 32214 59712 32220 59724
rect 32272 59712 32278 59764
rect 36538 59752 36544 59764
rect 36499 59724 36544 59752
rect 36538 59712 36544 59724
rect 36596 59712 36602 59764
rect 44082 59752 44088 59764
rect 44043 59724 44088 59752
rect 44082 59712 44088 59724
rect 44140 59712 44146 59764
rect 31754 59684 31760 59696
rect 27356 59656 31760 59684
rect 27218 59647 27276 59653
rect 31754 59644 31760 59656
rect 31812 59644 31818 59696
rect 33962 59684 33968 59696
rect 32508 59656 33824 59684
rect 33923 59656 33968 59684
rect 25225 59619 25283 59625
rect 25225 59585 25237 59619
rect 25271 59585 25283 59619
rect 25225 59579 25283 59585
rect 25317 59619 25375 59625
rect 25317 59585 25329 59619
rect 25363 59616 25375 59619
rect 25406 59616 25412 59628
rect 25363 59588 25412 59616
rect 25363 59585 25375 59588
rect 25317 59579 25375 59585
rect 25406 59576 25412 59588
rect 25464 59576 25470 59628
rect 26970 59616 26976 59628
rect 26931 59588 26976 59616
rect 26970 59576 26976 59588
rect 27028 59576 27034 59628
rect 27614 59576 27620 59628
rect 27672 59616 27678 59628
rect 28534 59616 28540 59628
rect 27672 59588 28540 59616
rect 27672 59576 27678 59588
rect 28534 59576 28540 59588
rect 28592 59616 28598 59628
rect 28902 59616 28908 59628
rect 28592 59588 28908 59616
rect 28592 59576 28598 59588
rect 28902 59576 28908 59588
rect 28960 59576 28966 59628
rect 29638 59625 29644 59628
rect 29632 59616 29644 59625
rect 29599 59588 29644 59616
rect 29632 59579 29644 59588
rect 29638 59576 29644 59579
rect 29696 59576 29702 59628
rect 32508 59625 32536 59656
rect 33796 59628 33824 59656
rect 33962 59644 33968 59656
rect 34020 59644 34026 59696
rect 35621 59687 35679 59693
rect 35621 59653 35633 59687
rect 35667 59684 35679 59687
rect 53834 59684 53840 59696
rect 35667 59656 53840 59684
rect 35667 59653 35679 59656
rect 35621 59647 35679 59653
rect 53834 59644 53840 59656
rect 53892 59644 53898 59696
rect 32493 59619 32551 59625
rect 32493 59585 32505 59619
rect 32539 59585 32551 59619
rect 32493 59579 32551 59585
rect 32585 59619 32643 59625
rect 32585 59585 32597 59619
rect 32631 59585 32643 59619
rect 32585 59579 32643 59585
rect 1854 59548 1860 59560
rect 1815 59520 1860 59548
rect 1854 59508 1860 59520
rect 1912 59508 1918 59560
rect 2774 59548 2780 59560
rect 2735 59520 2780 59548
rect 2774 59508 2780 59520
rect 2832 59508 2838 59560
rect 16669 59551 16727 59557
rect 16669 59517 16681 59551
rect 16715 59548 16727 59551
rect 16942 59548 16948 59560
rect 16715 59520 16948 59548
rect 16715 59517 16727 59520
rect 16669 59511 16727 59517
rect 16942 59508 16948 59520
rect 17000 59548 17006 59560
rect 19638 59551 19696 59557
rect 19638 59548 19650 59551
rect 17000 59520 19650 59548
rect 17000 59508 17006 59520
rect 19638 59517 19650 59520
rect 19684 59517 19696 59551
rect 19638 59511 19696 59517
rect 19797 59551 19855 59557
rect 19797 59517 19809 59551
rect 19843 59548 19855 59551
rect 19978 59548 19984 59560
rect 19843 59520 19984 59548
rect 19843 59517 19855 59520
rect 19797 59511 19855 59517
rect 19978 59508 19984 59520
rect 20036 59508 20042 59560
rect 29362 59548 29368 59560
rect 29323 59520 29368 59548
rect 29362 59508 29368 59520
rect 29420 59508 29426 59560
rect 31570 59508 31576 59560
rect 31628 59548 31634 59560
rect 32600 59548 32628 59579
rect 32674 59576 32680 59628
rect 32732 59616 32738 59628
rect 32732 59588 32777 59616
rect 32732 59576 32738 59588
rect 32858 59576 32864 59628
rect 32916 59616 32922 59628
rect 33778 59616 33784 59628
rect 32916 59588 32961 59616
rect 33739 59588 33784 59616
rect 32916 59576 32922 59588
rect 33778 59576 33784 59588
rect 33836 59576 33842 59628
rect 37366 59576 37372 59628
rect 37424 59616 37430 59628
rect 37533 59619 37591 59625
rect 37533 59616 37545 59619
rect 37424 59588 37545 59616
rect 37424 59576 37430 59588
rect 37533 59585 37545 59588
rect 37579 59585 37591 59619
rect 39666 59616 39672 59628
rect 39627 59588 39672 59616
rect 37533 59579 37591 59585
rect 39666 59576 39672 59588
rect 39724 59576 39730 59628
rect 41417 59619 41475 59625
rect 41417 59585 41429 59619
rect 41463 59585 41475 59619
rect 41598 59616 41604 59628
rect 41559 59588 41604 59616
rect 41417 59579 41475 59585
rect 31628 59520 32628 59548
rect 31628 59508 31634 59520
rect 35986 59508 35992 59560
rect 36044 59548 36050 59560
rect 36081 59551 36139 59557
rect 36081 59548 36093 59551
rect 36044 59520 36093 59548
rect 36044 59508 36050 59520
rect 36081 59517 36093 59520
rect 36127 59548 36139 59551
rect 36262 59548 36268 59560
rect 36127 59520 36268 59548
rect 36127 59517 36139 59520
rect 36081 59511 36139 59517
rect 36262 59508 36268 59520
rect 36320 59508 36326 59560
rect 37274 59548 37280 59560
rect 37235 59520 37280 59548
rect 37274 59508 37280 59520
rect 37332 59508 37338 59560
rect 39206 59508 39212 59560
rect 39264 59548 39270 59560
rect 39393 59551 39451 59557
rect 39393 59548 39405 59551
rect 39264 59520 39405 59548
rect 39264 59508 39270 59520
rect 39393 59517 39405 59520
rect 39439 59517 39451 59551
rect 41432 59548 41460 59579
rect 41598 59576 41604 59588
rect 41656 59576 41662 59628
rect 41690 59576 41696 59628
rect 41748 59616 41754 59628
rect 41748 59588 41793 59616
rect 41748 59576 41754 59588
rect 42978 59576 42984 59628
rect 43036 59616 43042 59628
rect 43349 59619 43407 59625
rect 43349 59616 43361 59619
rect 43036 59588 43361 59616
rect 43036 59576 43042 59588
rect 43349 59585 43361 59588
rect 43395 59585 43407 59619
rect 43349 59579 43407 59585
rect 43530 59576 43536 59628
rect 43588 59616 43594 59628
rect 43993 59619 44051 59625
rect 43993 59616 44005 59619
rect 43588 59588 44005 59616
rect 43588 59576 43594 59588
rect 43993 59585 44005 59588
rect 44039 59585 44051 59619
rect 44174 59616 44180 59628
rect 44135 59588 44180 59616
rect 43993 59579 44051 59585
rect 44174 59576 44180 59588
rect 44232 59576 44238 59628
rect 67266 59616 67272 59628
rect 67227 59588 67272 59616
rect 67266 59576 67272 59588
rect 67324 59576 67330 59628
rect 41506 59548 41512 59560
rect 41432 59520 41512 59548
rect 39393 59511 39451 59517
rect 41506 59508 41512 59520
rect 41564 59508 41570 59560
rect 41708 59548 41736 59576
rect 42610 59548 42616 59560
rect 41708 59520 42616 59548
rect 42610 59508 42616 59520
rect 42668 59548 42674 59560
rect 43165 59551 43223 59557
rect 43165 59548 43177 59551
rect 42668 59520 43177 59548
rect 42668 59508 42674 59520
rect 43165 59517 43177 59520
rect 43211 59517 43223 59551
rect 43165 59511 43223 59517
rect 43257 59551 43315 59557
rect 43257 59517 43269 59551
rect 43303 59517 43315 59551
rect 43257 59511 43315 59517
rect 43441 59551 43499 59557
rect 43441 59517 43453 59551
rect 43487 59517 43499 59551
rect 43441 59511 43499 59517
rect 19242 59480 19248 59492
rect 19203 59452 19248 59480
rect 19242 59440 19248 59452
rect 19300 59440 19306 59492
rect 20441 59483 20499 59489
rect 20441 59449 20453 59483
rect 20487 59480 20499 59483
rect 22186 59480 22192 59492
rect 20487 59452 22192 59480
rect 20487 59449 20499 59452
rect 20441 59443 20499 59449
rect 22186 59440 22192 59452
rect 22244 59440 22250 59492
rect 36354 59480 36360 59492
rect 36315 59452 36360 59480
rect 36354 59440 36360 59452
rect 36412 59480 36418 59492
rect 36630 59480 36636 59492
rect 36412 59452 36636 59480
rect 36412 59440 36418 59452
rect 36630 59440 36636 59452
rect 36688 59440 36694 59492
rect 42702 59440 42708 59492
rect 42760 59480 42766 59492
rect 43272 59480 43300 59511
rect 42760 59452 43300 59480
rect 42760 59440 42766 59452
rect 14366 59372 14372 59424
rect 14424 59412 14430 59424
rect 14461 59415 14519 59421
rect 14461 59412 14473 59415
rect 14424 59384 14473 59412
rect 14424 59372 14430 59384
rect 14461 59381 14473 59384
rect 14507 59381 14519 59415
rect 14461 59375 14519 59381
rect 18782 59372 18788 59424
rect 18840 59412 18846 59424
rect 20346 59412 20352 59424
rect 18840 59384 20352 59412
rect 18840 59372 18846 59384
rect 20346 59372 20352 59384
rect 20404 59372 20410 59424
rect 22002 59372 22008 59424
rect 22060 59412 22066 59424
rect 24213 59415 24271 59421
rect 24213 59412 24225 59415
rect 22060 59384 24225 59412
rect 22060 59372 22066 59384
rect 24213 59381 24225 59384
rect 24259 59381 24271 59415
rect 24213 59375 24271 59381
rect 29270 59372 29276 59424
rect 29328 59412 29334 59424
rect 30745 59415 30803 59421
rect 30745 59412 30757 59415
rect 29328 59384 30757 59412
rect 29328 59372 29334 59384
rect 30745 59381 30757 59384
rect 30791 59381 30803 59415
rect 30745 59375 30803 59381
rect 38657 59415 38715 59421
rect 38657 59381 38669 59415
rect 38703 59412 38715 59415
rect 39114 59412 39120 59424
rect 38703 59384 39120 59412
rect 38703 59381 38715 59384
rect 38657 59375 38715 59381
rect 39114 59372 39120 59384
rect 39172 59372 39178 59424
rect 41414 59372 41420 59424
rect 41472 59412 41478 59424
rect 42981 59415 43039 59421
rect 41472 59384 41517 59412
rect 41472 59372 41478 59384
rect 42981 59381 42993 59415
rect 43027 59412 43039 59415
rect 43070 59412 43076 59424
rect 43027 59384 43076 59412
rect 43027 59381 43039 59384
rect 42981 59375 43039 59381
rect 43070 59372 43076 59384
rect 43128 59372 43134 59424
rect 43162 59372 43168 59424
rect 43220 59412 43226 59424
rect 43456 59412 43484 59511
rect 43220 59384 43484 59412
rect 43220 59372 43226 59384
rect 67174 59372 67180 59424
rect 67232 59412 67238 59424
rect 67361 59415 67419 59421
rect 67361 59412 67373 59415
rect 67232 59384 67373 59412
rect 67232 59372 67238 59384
rect 67361 59381 67373 59384
rect 67407 59381 67419 59415
rect 67361 59375 67419 59381
rect 1104 59322 68816 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 34934 59322
rect 34986 59270 34998 59322
rect 35050 59270 35062 59322
rect 35114 59270 35126 59322
rect 35178 59270 35190 59322
rect 35242 59270 65654 59322
rect 65706 59270 65718 59322
rect 65770 59270 65782 59322
rect 65834 59270 65846 59322
rect 65898 59270 65910 59322
rect 65962 59270 68816 59322
rect 1104 59248 68816 59270
rect 1854 59168 1860 59220
rect 1912 59208 1918 59220
rect 2041 59211 2099 59217
rect 2041 59208 2053 59211
rect 1912 59180 2053 59208
rect 1912 59168 1918 59180
rect 2041 59177 2053 59180
rect 2087 59177 2099 59211
rect 2041 59171 2099 59177
rect 17405 59211 17463 59217
rect 17405 59177 17417 59211
rect 17451 59208 17463 59211
rect 17494 59208 17500 59220
rect 17451 59180 17500 59208
rect 17451 59177 17463 59180
rect 17405 59171 17463 59177
rect 17494 59168 17500 59180
rect 17552 59168 17558 59220
rect 29733 59211 29791 59217
rect 29733 59208 29745 59211
rect 22066 59180 29745 59208
rect 15470 59140 15476 59152
rect 15383 59112 15476 59140
rect 15470 59100 15476 59112
rect 15528 59140 15534 59152
rect 19518 59140 19524 59152
rect 15528 59112 19524 59140
rect 15528 59100 15534 59112
rect 19518 59100 19524 59112
rect 19576 59100 19582 59152
rect 1949 59007 2007 59013
rect 1949 58973 1961 59007
rect 1995 59004 2007 59007
rect 2038 59004 2044 59016
rect 1995 58976 2044 59004
rect 1995 58973 2007 58976
rect 1949 58967 2007 58973
rect 2038 58964 2044 58976
rect 2096 59004 2102 59016
rect 5994 59004 6000 59016
rect 2096 58976 6000 59004
rect 2096 58964 2102 58976
rect 5994 58964 6000 58976
rect 6052 58964 6058 59016
rect 14090 59004 14096 59016
rect 14051 58976 14096 59004
rect 14090 58964 14096 58976
rect 14148 58964 14154 59016
rect 14366 59013 14372 59016
rect 14360 59004 14372 59013
rect 14327 58976 14372 59004
rect 14360 58967 14372 58976
rect 14366 58964 14372 58967
rect 14424 58964 14430 59016
rect 17586 59004 17592 59016
rect 17547 58976 17592 59004
rect 17586 58964 17592 58976
rect 17644 58964 17650 59016
rect 19426 59004 19432 59016
rect 19387 58976 19432 59004
rect 19426 58964 19432 58976
rect 19484 58964 19490 59016
rect 20162 59004 20168 59016
rect 20123 58976 20168 59004
rect 20162 58964 20168 58976
rect 20220 58964 20226 59016
rect 21266 58964 21272 59016
rect 21324 59004 21330 59016
rect 21637 59007 21695 59013
rect 21637 59004 21649 59007
rect 21324 58976 21649 59004
rect 21324 58964 21330 58976
rect 21637 58973 21649 58976
rect 21683 58973 21695 59007
rect 21637 58967 21695 58973
rect 20438 58896 20444 58948
rect 20496 58936 20502 58948
rect 22066 58936 22094 59180
rect 29733 59177 29745 59180
rect 29779 59177 29791 59211
rect 29914 59208 29920 59220
rect 29875 59180 29920 59208
rect 29733 59171 29791 59177
rect 29914 59168 29920 59180
rect 29972 59168 29978 59220
rect 31481 59211 31539 59217
rect 31481 59177 31493 59211
rect 31527 59208 31539 59211
rect 32674 59208 32680 59220
rect 31527 59180 32680 59208
rect 31527 59177 31539 59180
rect 31481 59171 31539 59177
rect 32674 59168 32680 59180
rect 32732 59168 32738 59220
rect 36262 59208 36268 59220
rect 36223 59180 36268 59208
rect 36262 59168 36268 59180
rect 36320 59168 36326 59220
rect 39850 59208 39856 59220
rect 39811 59180 39856 59208
rect 39850 59168 39856 59180
rect 39908 59168 39914 59220
rect 41598 59168 41604 59220
rect 41656 59208 41662 59220
rect 42245 59211 42303 59217
rect 42245 59208 42257 59211
rect 41656 59180 42257 59208
rect 41656 59168 41662 59180
rect 42245 59177 42257 59180
rect 42291 59177 42303 59211
rect 42245 59171 42303 59177
rect 42981 59211 43039 59217
rect 42981 59177 42993 59211
rect 43027 59208 43039 59211
rect 44174 59208 44180 59220
rect 43027 59180 44180 59208
rect 43027 59177 43039 59180
rect 42981 59171 43039 59177
rect 38948 59112 39712 59140
rect 37274 59072 37280 59084
rect 37108 59044 37280 59072
rect 25409 59007 25467 59013
rect 25409 58973 25421 59007
rect 25455 59004 25467 59007
rect 25590 59004 25596 59016
rect 25455 58976 25596 59004
rect 25455 58973 25467 58976
rect 25409 58967 25467 58973
rect 25590 58964 25596 58976
rect 25648 58964 25654 59016
rect 31662 59004 31668 59016
rect 31623 58976 31668 59004
rect 31662 58964 31668 58976
rect 31720 58964 31726 59016
rect 31941 59007 31999 59013
rect 31941 58973 31953 59007
rect 31987 58973 31999 59007
rect 31941 58967 31999 58973
rect 34885 59007 34943 59013
rect 34885 58973 34897 59007
rect 34931 59004 34943 59007
rect 37108 59004 37136 59044
rect 37274 59032 37280 59044
rect 37332 59032 37338 59084
rect 38948 59081 38976 59112
rect 39684 59084 39712 59112
rect 38657 59075 38715 59081
rect 38657 59072 38669 59075
rect 37384 59044 38669 59072
rect 37384 59013 37412 59044
rect 38657 59041 38669 59044
rect 38703 59041 38715 59075
rect 38657 59035 38715 59041
rect 38933 59075 38991 59081
rect 38933 59041 38945 59075
rect 38979 59041 38991 59075
rect 39114 59072 39120 59084
rect 39075 59044 39120 59072
rect 38933 59035 38991 59041
rect 39114 59032 39120 59044
rect 39172 59032 39178 59084
rect 39666 59032 39672 59084
rect 39724 59072 39730 59084
rect 40129 59075 40187 59081
rect 40129 59072 40141 59075
rect 39724 59044 40141 59072
rect 39724 59032 39730 59044
rect 40129 59041 40141 59044
rect 40175 59041 40187 59075
rect 40129 59035 40187 59041
rect 40218 59032 40224 59084
rect 40276 59072 40282 59084
rect 40276 59044 40321 59072
rect 40276 59032 40282 59044
rect 34931 58976 37136 59004
rect 37185 59007 37243 59013
rect 34931 58973 34943 58976
rect 34885 58967 34943 58973
rect 37185 58973 37197 59007
rect 37231 58973 37243 59007
rect 37185 58967 37243 58973
rect 37369 59007 37427 59013
rect 37369 58973 37381 59007
rect 37415 58973 37427 59007
rect 38838 59004 38844 59016
rect 38799 58976 38844 59004
rect 37369 58967 37427 58973
rect 20496 58908 22094 58936
rect 20496 58896 20502 58908
rect 29270 58896 29276 58948
rect 29328 58936 29334 58948
rect 29549 58939 29607 58945
rect 29549 58936 29561 58939
rect 29328 58908 29561 58936
rect 29328 58896 29334 58908
rect 29549 58905 29561 58908
rect 29595 58905 29607 58939
rect 29549 58899 29607 58905
rect 30926 58896 30932 58948
rect 30984 58936 30990 58948
rect 31956 58936 31984 58967
rect 30984 58908 31984 58936
rect 35152 58939 35210 58945
rect 30984 58896 30990 58908
rect 35152 58905 35164 58939
rect 35198 58936 35210 58939
rect 35342 58936 35348 58948
rect 35198 58908 35348 58936
rect 35198 58905 35210 58908
rect 35152 58899 35210 58905
rect 35342 58896 35348 58908
rect 35400 58896 35406 58948
rect 37200 58936 37228 58967
rect 38838 58964 38844 58976
rect 38896 58964 38902 59016
rect 39025 59007 39083 59013
rect 39025 58973 39037 59007
rect 39071 58998 39083 59007
rect 39071 58973 39160 58998
rect 39025 58970 39160 58973
rect 39025 58967 39083 58970
rect 38010 58936 38016 58948
rect 37200 58908 38016 58936
rect 38010 58896 38016 58908
rect 38068 58896 38074 58948
rect 39132 58936 39160 58970
rect 39942 58964 39948 59016
rect 40000 59004 40006 59016
rect 40037 59007 40095 59013
rect 40037 59004 40049 59007
rect 40000 58976 40049 59004
rect 40000 58964 40006 58976
rect 40037 58973 40049 58976
rect 40083 58973 40095 59007
rect 40037 58967 40095 58973
rect 40310 58964 40316 59016
rect 40368 59004 40374 59016
rect 40368 58976 40413 59004
rect 40368 58964 40374 58976
rect 40770 58964 40776 59016
rect 40828 59004 40834 59016
rect 40865 59007 40923 59013
rect 40865 59004 40877 59007
rect 40828 58976 40877 59004
rect 40828 58964 40834 58976
rect 40865 58973 40877 58976
rect 40911 58973 40923 59007
rect 42260 59004 42288 59171
rect 44174 59168 44180 59180
rect 44232 59168 44238 59220
rect 42610 59032 42616 59084
rect 42668 59072 42674 59084
rect 42668 59044 43300 59072
rect 42668 59032 42674 59044
rect 42702 59004 42708 59016
rect 42260 58976 42708 59004
rect 40865 58967 40923 58973
rect 42702 58964 42708 58976
rect 42760 59004 42766 59016
rect 43272 59013 43300 59044
rect 43165 59007 43223 59013
rect 43165 59004 43177 59007
rect 42760 58976 43177 59004
rect 42760 58964 42766 58976
rect 43165 58973 43177 58976
rect 43211 58973 43223 59007
rect 43165 58967 43223 58973
rect 43257 59007 43315 59013
rect 43257 58973 43269 59007
rect 43303 59004 43315 59007
rect 43438 59004 43444 59016
rect 43303 58976 43444 59004
rect 43303 58973 43315 58976
rect 43257 58967 43315 58973
rect 43438 58964 43444 58976
rect 43496 58964 43502 59016
rect 40218 58936 40224 58948
rect 39132 58908 40224 58936
rect 40218 58896 40224 58908
rect 40276 58896 40282 58948
rect 41132 58939 41190 58945
rect 41132 58905 41144 58939
rect 41178 58936 41190 58939
rect 41230 58936 41236 58948
rect 41178 58908 41236 58936
rect 41178 58905 41190 58908
rect 41132 58899 41190 58905
rect 41230 58896 41236 58908
rect 41288 58896 41294 58948
rect 42978 58936 42984 58948
rect 42939 58908 42984 58936
rect 42978 58896 42984 58908
rect 43036 58896 43042 58948
rect 19058 58828 19064 58880
rect 19116 58868 19122 58880
rect 19429 58871 19487 58877
rect 19429 58868 19441 58871
rect 19116 58840 19441 58868
rect 19116 58828 19122 58840
rect 19429 58837 19441 58840
rect 19475 58837 19487 58871
rect 19978 58868 19984 58880
rect 19939 58840 19984 58868
rect 19429 58831 19487 58837
rect 19978 58828 19984 58840
rect 20036 58828 20042 58880
rect 21450 58868 21456 58880
rect 21411 58840 21456 58868
rect 21450 58828 21456 58840
rect 21508 58828 21514 58880
rect 25222 58868 25228 58880
rect 25183 58840 25228 58868
rect 25222 58828 25228 58840
rect 25280 58828 25286 58880
rect 29759 58871 29817 58877
rect 29759 58837 29771 58871
rect 29805 58868 29817 58871
rect 30466 58868 30472 58880
rect 29805 58840 30472 58868
rect 29805 58837 29817 58840
rect 29759 58831 29817 58837
rect 30466 58828 30472 58840
rect 30524 58828 30530 58880
rect 31754 58828 31760 58880
rect 31812 58868 31818 58880
rect 31849 58871 31907 58877
rect 31849 58868 31861 58871
rect 31812 58840 31861 58868
rect 31812 58828 31818 58840
rect 31849 58837 31861 58840
rect 31895 58837 31907 58871
rect 31849 58831 31907 58837
rect 37458 58828 37464 58880
rect 37516 58868 37522 58880
rect 37553 58871 37611 58877
rect 37553 58868 37565 58871
rect 37516 58840 37565 58868
rect 37516 58828 37522 58840
rect 37553 58837 37565 58840
rect 37599 58837 37611 58871
rect 37553 58831 37611 58837
rect 38838 58828 38844 58880
rect 38896 58868 38902 58880
rect 39942 58868 39948 58880
rect 38896 58840 39948 58868
rect 38896 58828 38902 58840
rect 39942 58828 39948 58840
rect 40000 58828 40006 58880
rect 1104 58778 68816 58800
rect 1104 58726 19574 58778
rect 19626 58726 19638 58778
rect 19690 58726 19702 58778
rect 19754 58726 19766 58778
rect 19818 58726 19830 58778
rect 19882 58726 50294 58778
rect 50346 58726 50358 58778
rect 50410 58726 50422 58778
rect 50474 58726 50486 58778
rect 50538 58726 50550 58778
rect 50602 58726 68816 58778
rect 1104 58704 68816 58726
rect 14090 58664 14096 58676
rect 14051 58636 14096 58664
rect 14090 58624 14096 58636
rect 14148 58624 14154 58676
rect 14642 58624 14648 58676
rect 14700 58664 14706 58676
rect 15105 58667 15163 58673
rect 15105 58664 15117 58667
rect 14700 58636 15117 58664
rect 14700 58624 14706 58636
rect 15105 58633 15117 58636
rect 15151 58633 15163 58667
rect 15105 58627 15163 58633
rect 20346 58624 20352 58676
rect 20404 58664 20410 58676
rect 20441 58667 20499 58673
rect 20441 58664 20453 58667
rect 20404 58636 20453 58664
rect 20404 58624 20410 58636
rect 20441 58633 20453 58636
rect 20487 58633 20499 58667
rect 20441 58627 20499 58633
rect 20622 58624 20628 58676
rect 20680 58664 20686 58676
rect 21101 58667 21159 58673
rect 21101 58664 21113 58667
rect 20680 58636 21113 58664
rect 20680 58624 20686 58636
rect 21101 58633 21113 58636
rect 21147 58633 21159 58667
rect 21266 58664 21272 58676
rect 21227 58636 21272 58664
rect 21101 58627 21159 58633
rect 21266 58624 21272 58636
rect 21324 58624 21330 58676
rect 23201 58667 23259 58673
rect 23201 58664 23213 58667
rect 21376 58636 23213 58664
rect 15470 58596 15476 58608
rect 14844 58568 15476 58596
rect 13814 58488 13820 58540
rect 13872 58528 13878 58540
rect 14844 58537 14872 58568
rect 15470 58556 15476 58568
rect 15528 58556 15534 58608
rect 19328 58599 19386 58605
rect 19328 58565 19340 58599
rect 19374 58596 19386 58599
rect 19978 58596 19984 58608
rect 19374 58568 19984 58596
rect 19374 58565 19386 58568
rect 19328 58559 19386 58565
rect 19978 58556 19984 58568
rect 20036 58556 20042 58608
rect 20901 58599 20959 58605
rect 20901 58565 20913 58599
rect 20947 58596 20959 58599
rect 20990 58596 20996 58608
rect 20947 58568 20996 58596
rect 20947 58565 20959 58568
rect 20901 58559 20959 58565
rect 20990 58556 20996 58568
rect 21048 58556 21054 58608
rect 13909 58531 13967 58537
rect 13909 58528 13921 58531
rect 13872 58500 13921 58528
rect 13872 58488 13878 58500
rect 13909 58497 13921 58500
rect 13955 58497 13967 58531
rect 13909 58491 13967 58497
rect 14829 58531 14887 58537
rect 14829 58497 14841 58531
rect 14875 58497 14887 58531
rect 14829 58491 14887 58497
rect 14921 58531 14979 58537
rect 14921 58497 14933 58531
rect 14967 58528 14979 58531
rect 15194 58528 15200 58540
rect 14967 58500 15200 58528
rect 14967 58497 14979 58500
rect 14921 58491 14979 58497
rect 15194 58488 15200 58500
rect 15252 58528 15258 58540
rect 16022 58528 16028 58540
rect 15252 58500 16028 58528
rect 15252 58488 15258 58500
rect 16022 58488 16028 58500
rect 16080 58488 16086 58540
rect 17126 58528 17132 58540
rect 17087 58500 17132 58528
rect 17126 58488 17132 58500
rect 17184 58488 17190 58540
rect 19058 58528 19064 58540
rect 19019 58500 19064 58528
rect 19058 58488 19064 58500
rect 19116 58488 19122 58540
rect 21008 58528 21036 58556
rect 21376 58528 21404 58636
rect 23201 58633 23213 58636
rect 23247 58633 23259 58667
rect 25590 58664 25596 58676
rect 25551 58636 25596 58664
rect 23201 58627 23259 58633
rect 25590 58624 25596 58636
rect 25648 58624 25654 58676
rect 26234 58624 26240 58676
rect 26292 58664 26298 58676
rect 28902 58664 28908 58676
rect 26292 58636 28908 58664
rect 26292 58624 26298 58636
rect 28902 58624 28908 58636
rect 28960 58624 28966 58676
rect 31754 58624 31760 58676
rect 31812 58664 31818 58676
rect 32493 58667 32551 58673
rect 32493 58664 32505 58667
rect 31812 58636 32505 58664
rect 31812 58624 31818 58636
rect 32493 58633 32505 58636
rect 32539 58633 32551 58667
rect 32493 58627 32551 58633
rect 37277 58667 37335 58673
rect 37277 58633 37289 58667
rect 37323 58664 37335 58667
rect 37366 58664 37372 58676
rect 37323 58636 37372 58664
rect 37323 58633 37335 58636
rect 37277 58627 37335 58633
rect 37366 58624 37372 58636
rect 37424 58624 37430 58676
rect 39666 58624 39672 58676
rect 39724 58664 39730 58676
rect 39945 58667 40003 58673
rect 39945 58664 39957 58667
rect 39724 58636 39957 58664
rect 39724 58624 39730 58636
rect 39945 58633 39957 58636
rect 39991 58633 40003 58667
rect 41230 58664 41236 58676
rect 41191 58636 41236 58664
rect 39945 58627 40003 58633
rect 41230 58624 41236 58636
rect 41288 58624 41294 58676
rect 43257 58667 43315 58673
rect 43257 58633 43269 58667
rect 43303 58664 43315 58667
rect 43303 58636 43944 58664
rect 43303 58633 43315 58636
rect 43257 58627 43315 58633
rect 21450 58556 21456 58608
rect 21508 58596 21514 58608
rect 22066 58599 22124 58605
rect 22066 58596 22078 58599
rect 21508 58568 22078 58596
rect 21508 58556 21514 58568
rect 22066 58565 22078 58568
rect 22112 58565 22124 58599
rect 26252 58596 26280 58624
rect 22066 58559 22124 58565
rect 25332 58568 26280 58596
rect 24302 58528 24308 58540
rect 21008 58500 21404 58528
rect 24263 58500 24308 58528
rect 24302 58488 24308 58500
rect 24360 58488 24366 58540
rect 25332 58537 25360 58568
rect 27798 58556 27804 58608
rect 27856 58596 27862 58608
rect 29733 58599 29791 58605
rect 27856 58568 28120 58596
rect 27856 58556 27862 58568
rect 25317 58531 25375 58537
rect 25317 58497 25329 58531
rect 25363 58497 25375 58531
rect 25317 58491 25375 58497
rect 25406 58488 25412 58540
rect 25464 58528 25470 58540
rect 26329 58531 26387 58537
rect 25464 58500 25509 58528
rect 25464 58488 25470 58500
rect 26329 58497 26341 58531
rect 26375 58528 26387 58531
rect 26418 58528 26424 58540
rect 26375 58500 26424 58528
rect 26375 58497 26387 58500
rect 26329 58491 26387 58497
rect 26418 58488 26424 58500
rect 26476 58488 26482 58540
rect 27341 58531 27399 58537
rect 27341 58497 27353 58531
rect 27387 58528 27399 58531
rect 27706 58528 27712 58540
rect 27387 58500 27712 58528
rect 27387 58497 27399 58500
rect 27341 58491 27399 58497
rect 27706 58488 27712 58500
rect 27764 58488 27770 58540
rect 27890 58528 27896 58540
rect 27851 58500 27896 58528
rect 27890 58488 27896 58500
rect 27948 58488 27954 58540
rect 28092 58528 28120 58568
rect 29733 58565 29745 58599
rect 29779 58596 29791 58599
rect 29779 58568 32628 58596
rect 29779 58565 29791 58568
rect 29733 58559 29791 58565
rect 28092 58500 28304 58528
rect 20990 58420 20996 58472
rect 21048 58460 21054 58472
rect 21821 58463 21879 58469
rect 21821 58460 21833 58463
rect 21048 58432 21833 58460
rect 21048 58420 21054 58432
rect 21821 58429 21833 58432
rect 21867 58429 21879 58463
rect 21821 58423 21879 58429
rect 28077 58463 28135 58469
rect 28077 58429 28089 58463
rect 28123 58429 28135 58463
rect 28276 58460 28304 58500
rect 28902 58488 28908 58540
rect 28960 58537 28966 58540
rect 28960 58531 28988 58537
rect 28976 58497 28988 58531
rect 29086 58528 29092 58540
rect 29047 58500 29092 58528
rect 28960 58491 28988 58497
rect 28960 58488 28966 58491
rect 29086 58488 29092 58500
rect 29144 58488 29150 58540
rect 29822 58488 29828 58540
rect 29880 58528 29886 58540
rect 30193 58531 30251 58537
rect 30193 58528 30205 58531
rect 29880 58500 30205 58528
rect 29880 58488 29886 58500
rect 30193 58497 30205 58500
rect 30239 58497 30251 58531
rect 31294 58528 31300 58540
rect 31255 58500 31300 58528
rect 30193 58491 30251 58497
rect 31294 58488 31300 58500
rect 31352 58488 31358 58540
rect 31662 58488 31668 58540
rect 31720 58528 31726 58540
rect 32600 58537 32628 58568
rect 35342 58556 35348 58608
rect 35400 58596 35406 58608
rect 38105 58599 38163 58605
rect 38105 58596 38117 58599
rect 35400 58568 38117 58596
rect 35400 58556 35406 58568
rect 38105 58565 38117 58568
rect 38151 58565 38163 58599
rect 38105 58559 38163 58565
rect 38289 58599 38347 58605
rect 38289 58565 38301 58599
rect 38335 58596 38347 58599
rect 38746 58596 38752 58608
rect 38335 58568 38752 58596
rect 38335 58565 38347 58568
rect 38289 58559 38347 58565
rect 38746 58556 38752 58568
rect 38804 58556 38810 58608
rect 39114 58596 39120 58608
rect 39040 58568 39120 58596
rect 32309 58531 32367 58537
rect 32309 58528 32321 58531
rect 31720 58500 32321 58528
rect 31720 58488 31726 58500
rect 32309 58497 32321 58500
rect 32355 58497 32367 58531
rect 32309 58491 32367 58497
rect 32585 58531 32643 58537
rect 32585 58497 32597 58531
rect 32631 58497 32643 58531
rect 32585 58491 32643 58497
rect 33597 58531 33655 58537
rect 33597 58497 33609 58531
rect 33643 58528 33655 58531
rect 33686 58528 33692 58540
rect 33643 58500 33692 58528
rect 33643 58497 33655 58500
rect 33597 58491 33655 58497
rect 33686 58488 33692 58500
rect 33744 58488 33750 58540
rect 37458 58528 37464 58540
rect 37419 58500 37464 58528
rect 37458 58488 37464 58500
rect 37516 58488 37522 58540
rect 39040 58537 39068 58568
rect 39114 58556 39120 58568
rect 39172 58556 39178 58608
rect 39761 58599 39819 58605
rect 39761 58565 39773 58599
rect 39807 58596 39819 58599
rect 41506 58596 41512 58608
rect 39807 58568 41512 58596
rect 39807 58565 39819 58568
rect 39761 58559 39819 58565
rect 41506 58556 41512 58568
rect 41564 58556 41570 58608
rect 39025 58531 39083 58537
rect 39025 58497 39037 58531
rect 39071 58497 39083 58531
rect 39206 58528 39212 58540
rect 39167 58500 39212 58528
rect 39025 58491 39083 58497
rect 39206 58488 39212 58500
rect 39264 58488 39270 58540
rect 39942 58488 39948 58540
rect 40000 58528 40006 58540
rect 40037 58531 40095 58537
rect 40037 58528 40049 58531
rect 40000 58500 40049 58528
rect 40000 58488 40006 58500
rect 40037 58497 40049 58500
rect 40083 58497 40095 58531
rect 40037 58491 40095 58497
rect 40310 58488 40316 58540
rect 40368 58528 40374 58540
rect 40497 58531 40555 58537
rect 40497 58528 40509 58531
rect 40368 58500 40509 58528
rect 40368 58488 40374 58500
rect 40497 58497 40509 58500
rect 40543 58497 40555 58531
rect 40497 58491 40555 58497
rect 28534 58460 28540 58472
rect 28276 58432 28540 58460
rect 28077 58423 28135 58429
rect 16758 58284 16764 58336
rect 16816 58324 16822 58336
rect 16945 58327 17003 58333
rect 16945 58324 16957 58327
rect 16816 58296 16957 58324
rect 16816 58284 16822 58296
rect 16945 58293 16957 58296
rect 16991 58293 17003 58327
rect 16945 58287 17003 58293
rect 20438 58284 20444 58336
rect 20496 58324 20502 58336
rect 21085 58327 21143 58333
rect 21085 58324 21097 58327
rect 20496 58296 21097 58324
rect 20496 58284 20502 58296
rect 21085 58293 21097 58296
rect 21131 58293 21143 58327
rect 21085 58287 21143 58293
rect 24397 58327 24455 58333
rect 24397 58293 24409 58327
rect 24443 58324 24455 58327
rect 24578 58324 24584 58336
rect 24443 58296 24584 58324
rect 24443 58293 24455 58296
rect 24397 58287 24455 58293
rect 24578 58284 24584 58296
rect 24636 58284 24642 58336
rect 26326 58324 26332 58336
rect 26287 58296 26332 58324
rect 26326 58284 26332 58296
rect 26384 58284 26390 58336
rect 26970 58284 26976 58336
rect 27028 58324 27034 58336
rect 27157 58327 27215 58333
rect 27157 58324 27169 58327
rect 27028 58296 27169 58324
rect 27028 58284 27034 58296
rect 27157 58293 27169 58296
rect 27203 58293 27215 58327
rect 28092 58324 28120 58423
rect 28534 58420 28540 58432
rect 28592 58420 28598 58472
rect 28810 58460 28816 58472
rect 28771 58432 28816 58460
rect 28810 58420 28816 58432
rect 28868 58420 28874 58472
rect 39301 58463 39359 58469
rect 39301 58429 39313 58463
rect 39347 58460 39359 58463
rect 40218 58460 40224 58472
rect 39347 58432 40224 58460
rect 39347 58429 39359 58432
rect 39301 58423 39359 58429
rect 40218 58420 40224 58432
rect 40276 58420 40282 58472
rect 40512 58460 40540 58491
rect 41414 58488 41420 58540
rect 41472 58528 41478 58540
rect 41472 58500 41517 58528
rect 41472 58488 41478 58500
rect 41598 58488 41604 58540
rect 41656 58528 41662 58540
rect 41693 58531 41751 58537
rect 41693 58528 41705 58531
rect 41656 58500 41705 58528
rect 41656 58488 41662 58500
rect 41693 58497 41705 58500
rect 41739 58497 41751 58531
rect 41693 58491 41751 58497
rect 42978 58488 42984 58540
rect 43036 58528 43042 58540
rect 43625 58531 43683 58537
rect 43036 58526 43576 58528
rect 43625 58526 43637 58531
rect 43036 58500 43637 58526
rect 43036 58488 43042 58500
rect 43548 58498 43637 58500
rect 43625 58497 43637 58498
rect 43671 58497 43683 58531
rect 43916 58528 43944 58636
rect 44453 58531 44511 58537
rect 44453 58528 44465 58531
rect 43916 58500 44465 58528
rect 43625 58491 43683 58497
rect 44453 58497 44465 58500
rect 44499 58497 44511 58531
rect 44453 58491 44511 58497
rect 43162 58460 43168 58472
rect 40512 58432 43168 58460
rect 43162 58420 43168 58432
rect 43220 58420 43226 58472
rect 43438 58460 43444 58472
rect 43399 58432 43444 58460
rect 43438 58420 43444 58432
rect 43496 58420 43502 58472
rect 43533 58463 43591 58469
rect 43533 58429 43545 58463
rect 43579 58429 43591 58463
rect 43533 58423 43591 58429
rect 38930 58352 38936 58404
rect 38988 58392 38994 58404
rect 39761 58395 39819 58401
rect 39761 58392 39773 58395
rect 38988 58364 39773 58392
rect 38988 58352 38994 58364
rect 39761 58361 39773 58364
rect 39807 58361 39819 58395
rect 39761 58355 39819 58361
rect 42702 58352 42708 58404
rect 42760 58392 42766 58404
rect 43548 58392 43576 58423
rect 43714 58420 43720 58472
rect 43772 58460 43778 58472
rect 43772 58432 43817 58460
rect 43772 58420 43778 58432
rect 43898 58420 43904 58472
rect 43956 58460 43962 58472
rect 44269 58463 44327 58469
rect 44269 58460 44281 58463
rect 43956 58432 44281 58460
rect 43956 58420 43962 58432
rect 44269 58429 44281 58432
rect 44315 58429 44327 58463
rect 44269 58423 44327 58429
rect 42760 58364 43576 58392
rect 42760 58352 42766 58364
rect 29914 58324 29920 58336
rect 28092 58296 29920 58324
rect 27157 58287 27215 58293
rect 29914 58284 29920 58296
rect 29972 58284 29978 58336
rect 30374 58324 30380 58336
rect 30335 58296 30380 58324
rect 30374 58284 30380 58296
rect 30432 58284 30438 58336
rect 31110 58324 31116 58336
rect 31071 58296 31116 58324
rect 31110 58284 31116 58296
rect 31168 58284 31174 58336
rect 32125 58327 32183 58333
rect 32125 58293 32137 58327
rect 32171 58324 32183 58327
rect 32582 58324 32588 58336
rect 32171 58296 32588 58324
rect 32171 58293 32183 58296
rect 32125 58287 32183 58293
rect 32582 58284 32588 58296
rect 32640 58284 32646 58336
rect 33689 58327 33747 58333
rect 33689 58293 33701 58327
rect 33735 58324 33747 58327
rect 33870 58324 33876 58336
rect 33735 58296 33876 58324
rect 33735 58293 33747 58296
rect 33689 58287 33747 58293
rect 33870 58284 33876 58296
rect 33928 58284 33934 58336
rect 38654 58284 38660 58336
rect 38712 58324 38718 58336
rect 38841 58327 38899 58333
rect 38841 58324 38853 58327
rect 38712 58296 38853 58324
rect 38712 58284 38718 58296
rect 38841 58293 38853 58296
rect 38887 58293 38899 58327
rect 38841 58287 38899 58293
rect 40681 58327 40739 58333
rect 40681 58293 40693 58327
rect 40727 58324 40739 58327
rect 41414 58324 41420 58336
rect 40727 58296 41420 58324
rect 40727 58293 40739 58296
rect 40681 58287 40739 58293
rect 41414 58284 41420 58296
rect 41472 58284 41478 58336
rect 41598 58324 41604 58336
rect 41559 58296 41604 58324
rect 41598 58284 41604 58296
rect 41656 58284 41662 58336
rect 44266 58284 44272 58336
rect 44324 58324 44330 58336
rect 44637 58327 44695 58333
rect 44637 58324 44649 58327
rect 44324 58296 44649 58324
rect 44324 58284 44330 58296
rect 44637 58293 44649 58296
rect 44683 58293 44695 58327
rect 44637 58287 44695 58293
rect 66254 58284 66260 58336
rect 66312 58324 66318 58336
rect 67637 58327 67695 58333
rect 67637 58324 67649 58327
rect 66312 58296 67649 58324
rect 66312 58284 66318 58296
rect 67637 58293 67649 58296
rect 67683 58293 67695 58327
rect 67637 58287 67695 58293
rect 1104 58234 68816 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 34934 58234
rect 34986 58182 34998 58234
rect 35050 58182 35062 58234
rect 35114 58182 35126 58234
rect 35178 58182 35190 58234
rect 35242 58182 65654 58234
rect 65706 58182 65718 58234
rect 65770 58182 65782 58234
rect 65834 58182 65846 58234
rect 65898 58182 65910 58234
rect 65962 58182 68816 58234
rect 1104 58160 68816 58182
rect 19981 58123 20039 58129
rect 19981 58089 19993 58123
rect 20027 58089 20039 58123
rect 20162 58120 20168 58132
rect 20123 58092 20168 58120
rect 19981 58083 20039 58089
rect 19996 58052 20024 58083
rect 20162 58080 20168 58092
rect 20220 58080 20226 58132
rect 20990 58120 20996 58132
rect 20951 58092 20996 58120
rect 20990 58080 20996 58092
rect 21048 58080 21054 58132
rect 28074 58120 28080 58132
rect 27987 58092 28080 58120
rect 28074 58080 28080 58092
rect 28132 58120 28138 58132
rect 28810 58120 28816 58132
rect 28132 58092 28816 58120
rect 28132 58080 28138 58092
rect 28810 58080 28816 58092
rect 28868 58080 28874 58132
rect 38010 58080 38016 58132
rect 38068 58120 38074 58132
rect 43898 58120 43904 58132
rect 38068 58092 43904 58120
rect 38068 58080 38074 58092
rect 43898 58080 43904 58092
rect 43956 58080 43962 58132
rect 20438 58052 20444 58064
rect 19996 58024 20444 58052
rect 20438 58012 20444 58024
rect 20496 58012 20502 58064
rect 38565 58055 38623 58061
rect 38565 58021 38577 58055
rect 38611 58052 38623 58055
rect 39022 58052 39028 58064
rect 38611 58024 39028 58052
rect 38611 58021 38623 58024
rect 38565 58015 38623 58021
rect 39022 58012 39028 58024
rect 39080 58012 39086 58064
rect 24578 57984 24584 57996
rect 24539 57956 24584 57984
rect 24578 57944 24584 57956
rect 24636 57944 24642 57996
rect 26142 57984 26148 57996
rect 26103 57956 26148 57984
rect 26142 57944 26148 57956
rect 26200 57944 26206 57996
rect 26326 57944 26332 57996
rect 26384 57984 26390 57996
rect 26697 57987 26755 57993
rect 26697 57984 26709 57987
rect 26384 57956 26709 57984
rect 26384 57944 26390 57956
rect 26697 57953 26709 57956
rect 26743 57953 26755 57987
rect 26697 57947 26755 57953
rect 15838 57916 15844 57928
rect 15799 57888 15844 57916
rect 15838 57876 15844 57888
rect 15896 57876 15902 57928
rect 16758 57925 16764 57928
rect 16025 57919 16083 57925
rect 16025 57885 16037 57919
rect 16071 57916 16083 57919
rect 16485 57919 16543 57925
rect 16485 57916 16497 57919
rect 16071 57888 16497 57916
rect 16071 57885 16083 57888
rect 16025 57879 16083 57885
rect 16485 57885 16497 57888
rect 16531 57885 16543 57919
rect 16752 57916 16764 57925
rect 16719 57888 16764 57916
rect 16485 57879 16543 57885
rect 16752 57879 16764 57888
rect 16758 57876 16764 57879
rect 16816 57876 16822 57928
rect 19426 57876 19432 57928
rect 19484 57916 19490 57928
rect 20809 57919 20867 57925
rect 20809 57916 20821 57919
rect 19484 57888 20821 57916
rect 19484 57876 19490 57888
rect 20809 57885 20821 57888
rect 20855 57885 20867 57919
rect 22462 57916 22468 57928
rect 22423 57888 22468 57916
rect 20809 57879 20867 57885
rect 22462 57876 22468 57888
rect 22520 57876 22526 57928
rect 26970 57925 26976 57928
rect 24397 57919 24455 57925
rect 24397 57916 24409 57919
rect 23860 57888 24409 57916
rect 19797 57851 19855 57857
rect 19797 57817 19809 57851
rect 19843 57848 19855 57851
rect 20346 57848 20352 57860
rect 19843 57820 20352 57848
rect 19843 57817 19855 57820
rect 19797 57811 19855 57817
rect 20346 57808 20352 57820
rect 20404 57808 20410 57860
rect 22738 57857 22744 57860
rect 22732 57811 22744 57857
rect 22796 57848 22802 57860
rect 22796 57820 22832 57848
rect 22738 57808 22744 57811
rect 22796 57808 22802 57820
rect 17862 57780 17868 57792
rect 17775 57752 17868 57780
rect 17862 57740 17868 57752
rect 17920 57780 17926 57792
rect 19150 57780 19156 57792
rect 17920 57752 19156 57780
rect 17920 57740 17926 57752
rect 19150 57740 19156 57752
rect 19208 57740 19214 57792
rect 19978 57740 19984 57792
rect 20036 57789 20042 57792
rect 20036 57783 20055 57789
rect 20043 57780 20055 57783
rect 20622 57780 20628 57792
rect 20043 57752 20628 57780
rect 20043 57749 20055 57752
rect 20036 57743 20055 57749
rect 20036 57740 20042 57743
rect 20622 57740 20628 57752
rect 20680 57740 20686 57792
rect 23014 57740 23020 57792
rect 23072 57780 23078 57792
rect 23860 57789 23888 57888
rect 24397 57885 24409 57888
rect 24443 57885 24455 57919
rect 26964 57916 26976 57925
rect 26931 57888 26976 57916
rect 24397 57879 24455 57885
rect 26964 57879 26976 57888
rect 26970 57876 26976 57879
rect 27028 57876 27034 57928
rect 29641 57919 29699 57925
rect 29641 57885 29653 57919
rect 29687 57916 29699 57919
rect 29822 57916 29828 57928
rect 29687 57888 29828 57916
rect 29687 57885 29699 57888
rect 29641 57879 29699 57885
rect 29822 57876 29828 57888
rect 29880 57876 29886 57928
rect 30285 57919 30343 57925
rect 30285 57885 30297 57919
rect 30331 57916 30343 57919
rect 30374 57916 30380 57928
rect 30331 57888 30380 57916
rect 30331 57885 30343 57888
rect 30285 57879 30343 57885
rect 30374 57876 30380 57888
rect 30432 57876 30438 57928
rect 30552 57919 30610 57925
rect 30552 57885 30564 57919
rect 30598 57916 30610 57919
rect 31110 57916 31116 57928
rect 30598 57888 31116 57916
rect 30598 57885 30610 57888
rect 30552 57879 30610 57885
rect 31110 57876 31116 57888
rect 31168 57876 31174 57928
rect 32401 57919 32459 57925
rect 32401 57885 32413 57919
rect 32447 57916 32459 57919
rect 33042 57916 33048 57928
rect 32447 57888 33048 57916
rect 32447 57885 32459 57888
rect 32401 57879 32459 57885
rect 33042 57876 33048 57888
rect 33100 57876 33106 57928
rect 34701 57919 34759 57925
rect 34701 57885 34713 57919
rect 34747 57916 34759 57919
rect 36262 57916 36268 57928
rect 34747 57888 36268 57916
rect 34747 57885 34759 57888
rect 34701 57879 34759 57885
rect 36262 57876 36268 57888
rect 36320 57876 36326 57928
rect 36909 57919 36967 57925
rect 36909 57885 36921 57919
rect 36955 57916 36967 57919
rect 37642 57916 37648 57928
rect 36955 57888 37648 57916
rect 36955 57885 36967 57888
rect 36909 57879 36967 57885
rect 37642 57876 37648 57888
rect 37700 57876 37706 57928
rect 38565 57919 38623 57925
rect 38565 57885 38577 57919
rect 38611 57916 38623 57919
rect 38654 57916 38660 57928
rect 38611 57888 38660 57916
rect 38611 57885 38623 57888
rect 38565 57879 38623 57885
rect 38654 57876 38660 57888
rect 38712 57876 38718 57928
rect 38749 57919 38807 57925
rect 38749 57885 38761 57919
rect 38795 57916 38807 57919
rect 38838 57916 38844 57928
rect 38795 57888 38844 57916
rect 38795 57885 38807 57888
rect 38749 57879 38807 57885
rect 38838 57876 38844 57888
rect 38896 57876 38902 57928
rect 44266 57916 44272 57928
rect 44227 57888 44272 57916
rect 44266 57876 44272 57888
rect 44324 57876 44330 57928
rect 45005 57919 45063 57925
rect 45005 57885 45017 57919
rect 45051 57885 45063 57919
rect 66254 57916 66260 57928
rect 66215 57888 66260 57916
rect 45005 57879 45063 57885
rect 29362 57808 29368 57860
rect 29420 57848 29426 57860
rect 29733 57851 29791 57857
rect 29733 57848 29745 57851
rect 29420 57820 29745 57848
rect 29420 57808 29426 57820
rect 29733 57817 29745 57820
rect 29779 57817 29791 57851
rect 29733 57811 29791 57817
rect 32122 57808 32128 57860
rect 32180 57848 32186 57860
rect 32646 57851 32704 57857
rect 32646 57848 32658 57851
rect 32180 57820 32658 57848
rect 32180 57808 32186 57820
rect 32646 57817 32658 57820
rect 32692 57817 32704 57851
rect 32646 57811 32704 57817
rect 33962 57808 33968 57860
rect 34020 57848 34026 57860
rect 34946 57851 35004 57857
rect 34946 57848 34958 57851
rect 34020 57820 34958 57848
rect 34020 57808 34026 57820
rect 34946 57817 34958 57820
rect 34992 57817 35004 57851
rect 34946 57811 35004 57817
rect 43070 57808 43076 57860
rect 43128 57848 43134 57860
rect 45020 57848 45048 57879
rect 66254 57876 66260 57888
rect 66312 57876 66318 57928
rect 68094 57916 68100 57928
rect 68055 57888 68100 57916
rect 68094 57876 68100 57888
rect 68152 57876 68158 57928
rect 45250 57851 45308 57857
rect 45250 57848 45262 57851
rect 43128 57820 45048 57848
rect 45112 57820 45262 57848
rect 43128 57808 43134 57820
rect 23845 57783 23903 57789
rect 23845 57780 23857 57783
rect 23072 57752 23857 57780
rect 23072 57740 23078 57752
rect 23845 57749 23857 57752
rect 23891 57749 23903 57783
rect 23845 57743 23903 57749
rect 29914 57740 29920 57792
rect 29972 57780 29978 57792
rect 31665 57783 31723 57789
rect 31665 57780 31677 57783
rect 29972 57752 31677 57780
rect 29972 57740 29978 57752
rect 31665 57749 31677 57752
rect 31711 57749 31723 57783
rect 31665 57743 31723 57749
rect 33686 57740 33692 57792
rect 33744 57780 33750 57792
rect 33781 57783 33839 57789
rect 33781 57780 33793 57783
rect 33744 57752 33793 57780
rect 33744 57740 33750 57752
rect 33781 57749 33793 57752
rect 33827 57749 33839 57783
rect 36078 57780 36084 57792
rect 36039 57752 36084 57780
rect 33781 57743 33839 57749
rect 36078 57740 36084 57752
rect 36136 57740 36142 57792
rect 36538 57740 36544 57792
rect 36596 57780 36602 57792
rect 36725 57783 36783 57789
rect 36725 57780 36737 57783
rect 36596 57752 36737 57780
rect 36596 57740 36602 57752
rect 36725 57749 36737 57752
rect 36771 57749 36783 57783
rect 36725 57743 36783 57749
rect 44085 57783 44143 57789
rect 44085 57749 44097 57783
rect 44131 57780 44143 57783
rect 45112 57780 45140 57820
rect 45250 57817 45262 57820
rect 45296 57817 45308 57851
rect 66438 57848 66444 57860
rect 66399 57820 66444 57848
rect 45250 57811 45308 57817
rect 66438 57808 66444 57820
rect 66496 57808 66502 57860
rect 46382 57780 46388 57792
rect 44131 57752 45140 57780
rect 46343 57752 46388 57780
rect 44131 57749 44143 57752
rect 44085 57743 44143 57749
rect 46382 57740 46388 57752
rect 46440 57740 46446 57792
rect 1104 57690 68816 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 68816 57690
rect 1104 57616 68816 57638
rect 17126 57536 17132 57588
rect 17184 57576 17190 57588
rect 17405 57579 17463 57585
rect 17405 57576 17417 57579
rect 17184 57548 17417 57576
rect 17184 57536 17190 57548
rect 17405 57545 17417 57548
rect 17451 57545 17463 57579
rect 19334 57576 19340 57588
rect 17405 57539 17463 57545
rect 18340 57548 19340 57576
rect 17862 57508 17868 57520
rect 17144 57480 17868 57508
rect 14636 57443 14694 57449
rect 14636 57409 14648 57443
rect 14682 57440 14694 57443
rect 14918 57440 14924 57452
rect 14682 57412 14924 57440
rect 14682 57409 14694 57412
rect 14636 57403 14694 57409
rect 14918 57400 14924 57412
rect 14976 57400 14982 57452
rect 17144 57449 17172 57480
rect 17862 57468 17868 57480
rect 17920 57468 17926 57520
rect 18340 57449 18368 57548
rect 19334 57536 19340 57548
rect 19392 57536 19398 57588
rect 22462 57536 22468 57588
rect 22520 57576 22526 57588
rect 30929 57579 30987 57585
rect 30929 57576 30941 57579
rect 22520 57548 30941 57576
rect 22520 57536 22526 57548
rect 30929 57545 30941 57548
rect 30975 57576 30987 57579
rect 33042 57576 33048 57588
rect 30975 57548 33048 57576
rect 30975 57545 30987 57548
rect 30929 57539 30987 57545
rect 33042 57536 33048 57548
rect 33100 57536 33106 57588
rect 36262 57536 36268 57588
rect 36320 57576 36326 57588
rect 37550 57576 37556 57588
rect 36320 57548 37556 57576
rect 36320 57536 36326 57548
rect 37550 57536 37556 57548
rect 37608 57576 37614 57588
rect 39669 57579 39727 57585
rect 39669 57576 39681 57579
rect 37608 57548 39681 57576
rect 37608 57536 37614 57548
rect 39669 57545 39681 57548
rect 39715 57576 39727 57579
rect 40770 57576 40776 57588
rect 39715 57548 40776 57576
rect 39715 57545 39727 57548
rect 39669 57539 39727 57545
rect 40770 57536 40776 57548
rect 40828 57536 40834 57588
rect 66438 57536 66444 57588
rect 66496 57576 66502 57588
rect 67545 57579 67603 57585
rect 67545 57576 67557 57579
rect 66496 57548 67557 57576
rect 66496 57536 66502 57548
rect 67545 57545 67557 57548
rect 67591 57545 67603 57579
rect 67545 57539 67603 57545
rect 22738 57508 22744 57520
rect 22699 57480 22744 57508
rect 22738 57468 22744 57480
rect 22796 57468 22802 57520
rect 25124 57511 25182 57517
rect 25124 57477 25136 57511
rect 25170 57508 25182 57511
rect 25222 57508 25228 57520
rect 25170 57480 25228 57508
rect 25170 57477 25182 57480
rect 25124 57471 25182 57477
rect 25222 57468 25228 57480
rect 25280 57468 25286 57520
rect 27706 57468 27712 57520
rect 27764 57508 27770 57520
rect 27801 57511 27859 57517
rect 27801 57508 27813 57511
rect 27764 57480 27813 57508
rect 27764 57468 27770 57480
rect 27801 57477 27813 57480
rect 27847 57477 27859 57511
rect 29914 57508 29920 57520
rect 29875 57480 29920 57508
rect 27801 57471 27859 57477
rect 29914 57468 29920 57480
rect 29972 57468 29978 57520
rect 30133 57511 30191 57517
rect 30133 57477 30145 57511
rect 30179 57508 30191 57511
rect 30466 57508 30472 57520
rect 30179 57480 30472 57508
rect 30179 57477 30191 57480
rect 30133 57471 30191 57477
rect 30466 57468 30472 57480
rect 30524 57468 30530 57520
rect 32122 57508 32128 57520
rect 32083 57480 32128 57508
rect 32122 57468 32128 57480
rect 32180 57468 32186 57520
rect 33870 57508 33876 57520
rect 32416 57480 33732 57508
rect 33831 57480 33876 57508
rect 17129 57443 17187 57449
rect 17129 57409 17141 57443
rect 17175 57409 17187 57443
rect 17129 57403 17187 57409
rect 17221 57443 17279 57449
rect 17221 57409 17233 57443
rect 17267 57409 17279 57443
rect 17221 57403 17279 57409
rect 18325 57443 18383 57449
rect 18325 57409 18337 57443
rect 18371 57409 18383 57443
rect 18325 57403 18383 57409
rect 14366 57372 14372 57384
rect 14327 57344 14372 57372
rect 14366 57332 14372 57344
rect 14424 57332 14430 57384
rect 16574 57332 16580 57384
rect 16632 57372 16638 57384
rect 17236 57372 17264 57403
rect 19150 57400 19156 57452
rect 19208 57449 19214 57452
rect 19208 57443 19236 57449
rect 19224 57409 19236 57443
rect 23014 57440 23020 57452
rect 22975 57412 23020 57440
rect 19208 57403 19236 57409
rect 19208 57400 19214 57403
rect 23014 57400 23020 57412
rect 23072 57400 23078 57452
rect 23109 57443 23167 57449
rect 23109 57409 23121 57443
rect 23155 57409 23167 57443
rect 23109 57403 23167 57409
rect 18138 57372 18144 57384
rect 16632 57344 17264 57372
rect 18099 57344 18144 57372
rect 16632 57332 16638 57344
rect 18138 57332 18144 57344
rect 18196 57332 18202 57384
rect 19061 57375 19119 57381
rect 19061 57372 19073 57375
rect 18432 57344 19073 57372
rect 15746 57304 15752 57316
rect 15659 57276 15752 57304
rect 15746 57264 15752 57276
rect 15804 57304 15810 57316
rect 18432 57304 18460 57344
rect 19061 57341 19073 57344
rect 19107 57341 19119 57375
rect 19061 57335 19119 57341
rect 19337 57375 19395 57381
rect 19337 57341 19349 57375
rect 19383 57372 19395 57375
rect 20070 57372 20076 57384
rect 19383 57344 20076 57372
rect 19383 57341 19395 57344
rect 19337 57335 19395 57341
rect 20070 57332 20076 57344
rect 20128 57332 20134 57384
rect 23124 57372 23152 57403
rect 23198 57400 23204 57452
rect 23256 57440 23262 57452
rect 23385 57443 23443 57449
rect 23256 57412 23301 57440
rect 23256 57400 23262 57412
rect 23385 57409 23397 57443
rect 23431 57440 23443 57443
rect 23658 57440 23664 57452
rect 23431 57412 23664 57440
rect 23431 57409 23443 57412
rect 23385 57403 23443 57409
rect 23658 57400 23664 57412
rect 23716 57400 23722 57452
rect 24305 57443 24363 57449
rect 24305 57409 24317 57443
rect 24351 57440 24363 57443
rect 24946 57440 24952 57452
rect 24351 57412 24952 57440
rect 24351 57409 24363 57412
rect 24305 57403 24363 57409
rect 24946 57400 24952 57412
rect 25004 57400 25010 57452
rect 27614 57440 27620 57452
rect 27575 57412 27620 57440
rect 27614 57400 27620 57412
rect 27672 57400 27678 57452
rect 30006 57400 30012 57452
rect 30064 57440 30070 57452
rect 32416 57449 32444 57480
rect 33704 57452 33732 57480
rect 33870 57468 33876 57480
rect 33928 57468 33934 57520
rect 37642 57508 37648 57520
rect 37603 57480 37648 57508
rect 37642 57468 37648 57480
rect 37700 57468 37706 57520
rect 38746 57468 38752 57520
rect 38804 57508 38810 57520
rect 39577 57511 39635 57517
rect 39577 57508 39589 57511
rect 38804 57480 39589 57508
rect 38804 57468 38810 57480
rect 39577 57477 39589 57480
rect 39623 57477 39635 57511
rect 39577 57471 39635 57477
rect 30837 57443 30895 57449
rect 30837 57440 30849 57443
rect 30064 57412 30849 57440
rect 30064 57400 30070 57412
rect 30837 57409 30849 57412
rect 30883 57409 30895 57443
rect 30837 57403 30895 57409
rect 32401 57443 32459 57449
rect 32401 57409 32413 57443
rect 32447 57409 32459 57443
rect 32401 57403 32459 57409
rect 32493 57443 32551 57449
rect 32493 57409 32505 57443
rect 32539 57409 32551 57443
rect 32493 57403 32551 57409
rect 24210 57372 24216 57384
rect 23124 57344 24216 57372
rect 24210 57332 24216 57344
rect 24268 57332 24274 57384
rect 24397 57375 24455 57381
rect 24397 57341 24409 57375
rect 24443 57372 24455 57375
rect 24857 57375 24915 57381
rect 24857 57372 24869 57375
rect 24443 57344 24869 57372
rect 24443 57341 24455 57344
rect 24397 57335 24455 57341
rect 24857 57341 24869 57344
rect 24903 57341 24915 57375
rect 24857 57335 24915 57341
rect 27433 57375 27491 57381
rect 27433 57341 27445 57375
rect 27479 57372 27491 57375
rect 28074 57372 28080 57384
rect 27479 57344 28080 57372
rect 27479 57341 27491 57344
rect 27433 57335 27491 57341
rect 28074 57332 28080 57344
rect 28132 57332 28138 57384
rect 30374 57332 30380 57384
rect 30432 57372 30438 57384
rect 31570 57372 31576 57384
rect 30432 57344 31576 57372
rect 30432 57332 30438 57344
rect 31570 57332 31576 57344
rect 31628 57372 31634 57384
rect 32508 57372 32536 57403
rect 32582 57400 32588 57452
rect 32640 57440 32646 57452
rect 32769 57443 32827 57449
rect 32640 57412 32685 57440
rect 32640 57400 32646 57412
rect 32769 57409 32781 57443
rect 32815 57440 32827 57443
rect 32858 57440 32864 57452
rect 32815 57412 32864 57440
rect 32815 57409 32827 57412
rect 32769 57403 32827 57409
rect 32858 57400 32864 57412
rect 32916 57440 32922 57452
rect 33686 57440 33692 57452
rect 32916 57412 33548 57440
rect 33647 57412 33692 57440
rect 32916 57400 32922 57412
rect 31628 57344 32536 57372
rect 31628 57332 31634 57344
rect 15804 57276 18460 57304
rect 18785 57307 18843 57313
rect 15804 57264 15810 57276
rect 18785 57273 18797 57307
rect 18831 57273 18843 57307
rect 26234 57304 26240 57316
rect 26195 57276 26240 57304
rect 18785 57267 18843 57273
rect 17954 57196 17960 57248
rect 18012 57236 18018 57248
rect 18800 57236 18828 57267
rect 26234 57264 26240 57276
rect 26292 57264 26298 57316
rect 30285 57307 30343 57313
rect 30285 57273 30297 57307
rect 30331 57304 30343 57307
rect 31294 57304 31300 57316
rect 30331 57276 31300 57304
rect 30331 57273 30343 57276
rect 30285 57267 30343 57273
rect 31294 57264 31300 57276
rect 31352 57264 31358 57316
rect 33520 57304 33548 57412
rect 33686 57400 33692 57412
rect 33744 57400 33750 57452
rect 36078 57440 36084 57452
rect 36039 57412 36084 57440
rect 36078 57400 36084 57412
rect 36136 57400 36142 57452
rect 36173 57443 36231 57449
rect 36173 57409 36185 57443
rect 36219 57440 36231 57443
rect 37366 57440 37372 57452
rect 36219 57412 37372 57440
rect 36219 57409 36231 57412
rect 36173 57403 36231 57409
rect 37366 57400 37372 57412
rect 37424 57440 37430 57452
rect 37461 57443 37519 57449
rect 37461 57440 37473 57443
rect 37424 57412 37473 57440
rect 37424 57400 37430 57412
rect 37461 57409 37473 57412
rect 37507 57409 37519 57443
rect 38838 57440 38844 57452
rect 37461 57403 37519 57409
rect 38120 57412 38844 57440
rect 34514 57372 34520 57384
rect 34475 57344 34520 57372
rect 34514 57332 34520 57344
rect 34572 57332 34578 57384
rect 37277 57375 37335 57381
rect 37277 57341 37289 57375
rect 37323 57372 37335 57375
rect 37642 57372 37648 57384
rect 37323 57344 37648 57372
rect 37323 57341 37335 57344
rect 37277 57335 37335 57341
rect 37642 57332 37648 57344
rect 37700 57372 37706 57384
rect 38120 57372 38148 57412
rect 38838 57400 38844 57412
rect 38896 57400 38902 57452
rect 41322 57440 41328 57452
rect 41283 57412 41328 57440
rect 41322 57400 41328 57412
rect 41380 57400 41386 57452
rect 42705 57443 42763 57449
rect 42705 57409 42717 57443
rect 42751 57440 42763 57443
rect 42978 57440 42984 57452
rect 42751 57412 42984 57440
rect 42751 57409 42763 57412
rect 42705 57403 42763 57409
rect 42978 57400 42984 57412
rect 43036 57440 43042 57452
rect 43714 57440 43720 57452
rect 43036 57412 43720 57440
rect 43036 57400 43042 57412
rect 43714 57400 43720 57412
rect 43772 57440 43778 57452
rect 46382 57440 46388 57452
rect 43772 57412 46388 57440
rect 43772 57400 43778 57412
rect 46382 57400 46388 57412
rect 46440 57400 46446 57452
rect 53098 57400 53104 57452
rect 53156 57440 53162 57452
rect 66990 57440 66996 57452
rect 53156 57412 66996 57440
rect 53156 57400 53162 57412
rect 66990 57400 66996 57412
rect 67048 57440 67054 57452
rect 67453 57443 67511 57449
rect 67453 57440 67465 57443
rect 67048 57412 67465 57440
rect 67048 57400 67054 57412
rect 67453 57409 67465 57412
rect 67499 57409 67511 57443
rect 67453 57403 67511 57409
rect 37700 57344 38148 57372
rect 37700 57332 37706 57344
rect 38654 57332 38660 57384
rect 38712 57372 38718 57384
rect 38749 57375 38807 57381
rect 38749 57372 38761 57375
rect 38712 57344 38761 57372
rect 38712 57332 38718 57344
rect 38749 57341 38761 57344
rect 38795 57341 38807 57375
rect 38749 57335 38807 57341
rect 38933 57375 38991 57381
rect 38933 57341 38945 57375
rect 38979 57372 38991 57375
rect 39114 57372 39120 57384
rect 38979 57344 39120 57372
rect 38979 57341 38991 57344
rect 38933 57335 38991 57341
rect 39114 57332 39120 57344
rect 39172 57332 39178 57384
rect 42794 57372 42800 57384
rect 42755 57344 42800 57372
rect 42794 57332 42800 57344
rect 42852 57332 42858 57384
rect 42886 57332 42892 57384
rect 42944 57372 42950 57384
rect 42944 57344 42989 57372
rect 42944 57332 42950 57344
rect 35894 57304 35900 57316
rect 33520 57276 35900 57304
rect 35894 57264 35900 57276
rect 35952 57304 35958 57316
rect 36170 57304 36176 57316
rect 35952 57276 36176 57304
rect 35952 57264 35958 57276
rect 36170 57264 36176 57276
rect 36228 57264 36234 57316
rect 19242 57236 19248 57248
rect 18012 57208 19248 57236
rect 18012 57196 18018 57208
rect 19242 57196 19248 57208
rect 19300 57196 19306 57248
rect 19981 57239 20039 57245
rect 19981 57205 19993 57239
rect 20027 57236 20039 57239
rect 22370 57236 22376 57248
rect 20027 57208 22376 57236
rect 20027 57205 20039 57208
rect 19981 57199 20039 57205
rect 22370 57196 22376 57208
rect 22428 57196 22434 57248
rect 30101 57239 30159 57245
rect 30101 57205 30113 57239
rect 30147 57236 30159 57239
rect 30190 57236 30196 57248
rect 30147 57208 30196 57236
rect 30147 57205 30159 57208
rect 30101 57199 30159 57205
rect 30190 57196 30196 57208
rect 30248 57196 30254 57248
rect 34146 57196 34152 57248
rect 34204 57236 34210 57248
rect 36357 57239 36415 57245
rect 36357 57236 36369 57239
rect 34204 57208 36369 57236
rect 34204 57196 34210 57208
rect 36357 57205 36369 57208
rect 36403 57205 36415 57239
rect 36357 57199 36415 57205
rect 38565 57239 38623 57245
rect 38565 57205 38577 57239
rect 38611 57236 38623 57239
rect 38930 57236 38936 57248
rect 38611 57208 38936 57236
rect 38611 57205 38623 57208
rect 38565 57199 38623 57205
rect 38930 57196 38936 57208
rect 38988 57196 38994 57248
rect 41138 57236 41144 57248
rect 41099 57208 41144 57236
rect 41138 57196 41144 57208
rect 41196 57196 41202 57248
rect 42521 57239 42579 57245
rect 42521 57205 42533 57239
rect 42567 57236 42579 57239
rect 42610 57236 42616 57248
rect 42567 57208 42616 57236
rect 42567 57205 42579 57208
rect 42521 57199 42579 57205
rect 42610 57196 42616 57208
rect 42668 57196 42674 57248
rect 1104 57146 68816 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 65654 57146
rect 65706 57094 65718 57146
rect 65770 57094 65782 57146
rect 65834 57094 65846 57146
rect 65898 57094 65910 57146
rect 65962 57094 68816 57146
rect 1104 57072 68816 57094
rect 14366 57032 14372 57044
rect 14327 57004 14372 57032
rect 14366 56992 14372 57004
rect 14424 56992 14430 57044
rect 21637 57035 21695 57041
rect 21637 57001 21649 57035
rect 21683 57032 21695 57035
rect 23198 57032 23204 57044
rect 21683 57004 23204 57032
rect 21683 57001 21695 57004
rect 21637 56995 21695 57001
rect 23198 56992 23204 57004
rect 23256 56992 23262 57044
rect 24210 56992 24216 57044
rect 24268 57032 24274 57044
rect 24949 57035 25007 57041
rect 24949 57032 24961 57035
rect 24268 57004 24961 57032
rect 24268 56992 24274 57004
rect 24949 57001 24961 57004
rect 24995 57032 25007 57035
rect 28169 57035 28227 57041
rect 24995 57004 28120 57032
rect 24995 57001 25007 57004
rect 24949 56995 25007 57001
rect 28092 56964 28120 57004
rect 28169 57001 28181 57035
rect 28215 57032 28227 57035
rect 28718 57032 28724 57044
rect 28215 57004 28724 57032
rect 28215 57001 28227 57004
rect 28169 56995 28227 57001
rect 28718 56992 28724 57004
rect 28776 56992 28782 57044
rect 33962 57032 33968 57044
rect 33923 57004 33968 57032
rect 33962 56992 33968 57004
rect 34020 56992 34026 57044
rect 37642 57032 37648 57044
rect 37603 57004 37648 57032
rect 37642 56992 37648 57004
rect 37700 56992 37706 57044
rect 38838 56992 38844 57044
rect 38896 57032 38902 57044
rect 39117 57035 39175 57041
rect 39117 57032 39129 57035
rect 38896 57004 39129 57032
rect 38896 56992 38902 57004
rect 39117 57001 39129 57004
rect 39163 57001 39175 57035
rect 39117 56995 39175 57001
rect 42886 56992 42892 57044
rect 42944 57032 42950 57044
rect 44453 57035 44511 57041
rect 44453 57032 44465 57035
rect 42944 57004 44465 57032
rect 42944 56992 42950 57004
rect 44453 57001 44465 57004
rect 44499 57001 44511 57035
rect 44453 56995 44511 57001
rect 30374 56964 30380 56976
rect 28092 56936 30380 56964
rect 30374 56924 30380 56936
rect 30432 56924 30438 56976
rect 34790 56924 34796 56976
rect 34848 56964 34854 56976
rect 35342 56964 35348 56976
rect 34848 56936 35348 56964
rect 34848 56924 34854 56936
rect 35342 56924 35348 56936
rect 35400 56924 35406 56976
rect 15013 56899 15071 56905
rect 15013 56865 15025 56899
rect 15059 56896 15071 56899
rect 15746 56896 15752 56908
rect 15059 56868 15752 56896
rect 15059 56865 15071 56868
rect 15013 56859 15071 56865
rect 15746 56856 15752 56868
rect 15804 56856 15810 56908
rect 18417 56899 18475 56905
rect 18417 56896 18429 56899
rect 17144 56868 18429 56896
rect 1394 56828 1400 56840
rect 1355 56800 1400 56828
rect 1394 56788 1400 56800
rect 1452 56788 1458 56840
rect 13814 56788 13820 56840
rect 13872 56828 13878 56840
rect 14185 56831 14243 56837
rect 14185 56828 14197 56831
rect 13872 56800 14197 56828
rect 13872 56788 13878 56800
rect 14185 56797 14197 56800
rect 14231 56797 14243 56831
rect 15194 56828 15200 56840
rect 15155 56800 15200 56828
rect 14185 56791 14243 56797
rect 15194 56788 15200 56800
rect 15252 56788 15258 56840
rect 17144 56837 17172 56868
rect 18417 56865 18429 56868
rect 18463 56865 18475 56899
rect 36262 56896 36268 56908
rect 36223 56868 36268 56896
rect 18417 56859 18475 56865
rect 36262 56856 36268 56868
rect 36320 56856 36326 56908
rect 40770 56896 40776 56908
rect 40731 56868 40776 56896
rect 40770 56856 40776 56868
rect 40828 56856 40834 56908
rect 43070 56896 43076 56908
rect 43031 56868 43076 56896
rect 43070 56856 43076 56868
rect 43128 56856 43134 56908
rect 17129 56831 17187 56837
rect 17129 56797 17141 56831
rect 17175 56797 17187 56831
rect 18138 56828 18144 56840
rect 18099 56800 18144 56828
rect 17129 56791 17187 56797
rect 18138 56788 18144 56800
rect 18196 56788 18202 56840
rect 18230 56788 18236 56840
rect 18288 56828 18294 56840
rect 18288 56800 18333 56828
rect 18288 56788 18294 56800
rect 19426 56788 19432 56840
rect 19484 56828 19490 56840
rect 19613 56831 19671 56837
rect 19613 56828 19625 56831
rect 19484 56800 19625 56828
rect 19484 56788 19490 56800
rect 19613 56797 19625 56800
rect 19659 56828 19671 56831
rect 19978 56828 19984 56840
rect 19659 56800 19984 56828
rect 19659 56797 19671 56800
rect 19613 56791 19671 56797
rect 19978 56788 19984 56800
rect 20036 56788 20042 56840
rect 20530 56828 20536 56840
rect 20491 56800 20536 56828
rect 20530 56788 20536 56800
rect 20588 56788 20594 56840
rect 21726 56788 21732 56840
rect 21784 56828 21790 56840
rect 21821 56831 21879 56837
rect 21821 56828 21833 56831
rect 21784 56800 21833 56828
rect 21784 56788 21790 56800
rect 21821 56797 21833 56800
rect 21867 56797 21879 56831
rect 21821 56791 21879 56797
rect 22097 56831 22155 56837
rect 22097 56797 22109 56831
rect 22143 56828 22155 56831
rect 22186 56828 22192 56840
rect 22143 56800 22192 56828
rect 22143 56797 22155 56800
rect 22097 56791 22155 56797
rect 22186 56788 22192 56800
rect 22244 56788 22250 56840
rect 26142 56828 26148 56840
rect 26103 56800 26148 56828
rect 26142 56788 26148 56800
rect 26200 56788 26206 56840
rect 30834 56828 30840 56840
rect 30795 56800 30840 56828
rect 30834 56788 30840 56800
rect 30892 56788 30898 56840
rect 33505 56831 33563 56837
rect 33505 56797 33517 56831
rect 33551 56797 33563 56831
rect 34146 56828 34152 56840
rect 34107 56800 34152 56828
rect 33505 56791 33563 56797
rect 24857 56763 24915 56769
rect 24857 56729 24869 56763
rect 24903 56760 24915 56763
rect 25038 56760 25044 56772
rect 24903 56732 25044 56760
rect 24903 56729 24915 56732
rect 24857 56723 24915 56729
rect 25038 56720 25044 56732
rect 25096 56720 25102 56772
rect 26412 56763 26470 56769
rect 26412 56729 26424 56763
rect 26458 56760 26470 56763
rect 26510 56760 26516 56772
rect 26458 56732 26516 56760
rect 26458 56729 26470 56732
rect 26412 56723 26470 56729
rect 26510 56720 26516 56732
rect 26568 56720 26574 56772
rect 28077 56763 28135 56769
rect 28077 56729 28089 56763
rect 28123 56760 28135 56763
rect 28626 56760 28632 56772
rect 28123 56732 28632 56760
rect 28123 56729 28135 56732
rect 28077 56723 28135 56729
rect 28626 56720 28632 56732
rect 28684 56720 28690 56772
rect 31104 56763 31162 56769
rect 31104 56729 31116 56763
rect 31150 56760 31162 56763
rect 31386 56760 31392 56772
rect 31150 56732 31392 56760
rect 31150 56729 31162 56732
rect 31104 56723 31162 56729
rect 31386 56720 31392 56732
rect 31444 56720 31450 56772
rect 33520 56760 33548 56791
rect 34146 56788 34152 56800
rect 34204 56788 34210 56840
rect 36538 56837 36544 56840
rect 36532 56828 36544 56837
rect 36499 56800 36544 56828
rect 36532 56791 36544 56800
rect 36538 56788 36544 56791
rect 36596 56788 36602 56840
rect 38930 56828 38936 56840
rect 38891 56800 38936 56828
rect 38930 56788 38936 56800
rect 38988 56788 38994 56840
rect 40788 56828 40816 56856
rect 42518 56828 42524 56840
rect 40788 56800 42524 56828
rect 42518 56788 42524 56800
rect 42576 56828 42582 56840
rect 43088 56828 43116 56856
rect 45370 56828 45376 56840
rect 42576 56800 43116 56828
rect 45331 56800 45376 56828
rect 42576 56788 42582 56800
rect 45370 56788 45376 56800
rect 45428 56788 45434 56840
rect 46842 56828 46848 56840
rect 46803 56800 46848 56828
rect 46842 56788 46848 56800
rect 46900 56788 46906 56840
rect 50341 56831 50399 56837
rect 50341 56797 50353 56831
rect 50387 56828 50399 56831
rect 50614 56828 50620 56840
rect 50387 56800 50620 56828
rect 50387 56797 50399 56800
rect 50341 56791 50399 56797
rect 50614 56788 50620 56800
rect 50672 56788 50678 56840
rect 67542 56788 67548 56840
rect 67600 56828 67606 56840
rect 67637 56831 67695 56837
rect 67637 56828 67649 56831
rect 67600 56800 67649 56828
rect 67600 56788 67606 56800
rect 67637 56797 67649 56800
rect 67683 56797 67695 56831
rect 67637 56791 67695 56797
rect 35066 56760 35072 56772
rect 33520 56732 35072 56760
rect 35066 56720 35072 56732
rect 35124 56720 35130 56772
rect 35161 56763 35219 56769
rect 35161 56729 35173 56763
rect 35207 56760 35219 56763
rect 35342 56760 35348 56772
rect 35207 56732 35348 56760
rect 35207 56729 35219 56732
rect 35161 56723 35219 56729
rect 35342 56720 35348 56732
rect 35400 56720 35406 56772
rect 38194 56720 38200 56772
rect 38252 56760 38258 56772
rect 38565 56763 38623 56769
rect 38565 56760 38577 56763
rect 38252 56732 38577 56760
rect 38252 56720 38258 56732
rect 38565 56729 38577 56732
rect 38611 56729 38623 56763
rect 38565 56723 38623 56729
rect 41040 56763 41098 56769
rect 41040 56729 41052 56763
rect 41086 56760 41098 56763
rect 41138 56760 41144 56772
rect 41086 56732 41144 56760
rect 41086 56729 41098 56732
rect 41040 56723 41098 56729
rect 41138 56720 41144 56732
rect 41196 56720 41202 56772
rect 43346 56769 43352 56772
rect 43340 56723 43352 56769
rect 43404 56760 43410 56772
rect 47112 56763 47170 56769
rect 43404 56732 43440 56760
rect 43346 56720 43352 56723
rect 43404 56720 43410 56732
rect 47112 56729 47124 56763
rect 47158 56760 47170 56763
rect 47578 56760 47584 56772
rect 47158 56732 47584 56760
rect 47158 56729 47170 56732
rect 47112 56723 47170 56729
rect 47578 56720 47584 56732
rect 47636 56720 47642 56772
rect 67913 56763 67971 56769
rect 67913 56760 67925 56763
rect 67284 56732 67925 56760
rect 1486 56652 1492 56704
rect 1544 56692 1550 56704
rect 1581 56695 1639 56701
rect 1581 56692 1593 56695
rect 1544 56664 1593 56692
rect 1544 56652 1550 56664
rect 1581 56661 1593 56664
rect 1627 56661 1639 56695
rect 15378 56692 15384 56704
rect 15339 56664 15384 56692
rect 1581 56655 1639 56661
rect 15378 56652 15384 56664
rect 15436 56652 15442 56704
rect 16942 56692 16948 56704
rect 16903 56664 16948 56692
rect 16942 56652 16948 56664
rect 17000 56652 17006 56704
rect 19426 56652 19432 56704
rect 19484 56692 19490 56704
rect 19797 56695 19855 56701
rect 19797 56692 19809 56695
rect 19484 56664 19809 56692
rect 19484 56652 19490 56664
rect 19797 56661 19809 56664
rect 19843 56661 19855 56695
rect 20346 56692 20352 56704
rect 20307 56664 20352 56692
rect 19797 56655 19855 56661
rect 20346 56652 20352 56664
rect 20404 56652 20410 56704
rect 22005 56695 22063 56701
rect 22005 56661 22017 56695
rect 22051 56692 22063 56695
rect 22186 56692 22192 56704
rect 22051 56664 22192 56692
rect 22051 56661 22063 56664
rect 22005 56655 22063 56661
rect 22186 56652 22192 56664
rect 22244 56652 22250 56704
rect 27522 56692 27528 56704
rect 27483 56664 27528 56692
rect 27522 56652 27528 56664
rect 27580 56652 27586 56704
rect 30374 56652 30380 56704
rect 30432 56692 30438 56704
rect 32217 56695 32275 56701
rect 32217 56692 32229 56695
rect 30432 56664 32229 56692
rect 30432 56652 30438 56664
rect 32217 56661 32229 56664
rect 32263 56661 32275 56695
rect 33318 56692 33324 56704
rect 33279 56664 33324 56692
rect 32217 56655 32275 56661
rect 33318 56652 33324 56664
rect 33376 56652 33382 56704
rect 38746 56692 38752 56704
rect 38707 56664 38752 56692
rect 38746 56652 38752 56664
rect 38804 56652 38810 56704
rect 38838 56652 38844 56704
rect 38896 56692 38902 56704
rect 38896 56664 38941 56692
rect 38896 56652 38902 56664
rect 40494 56652 40500 56704
rect 40552 56692 40558 56704
rect 42150 56692 42156 56704
rect 40552 56664 42156 56692
rect 40552 56652 40558 56664
rect 42150 56652 42156 56664
rect 42208 56652 42214 56704
rect 45186 56652 45192 56704
rect 45244 56692 45250 56704
rect 45373 56695 45431 56701
rect 45373 56692 45385 56695
rect 45244 56664 45385 56692
rect 45244 56652 45250 56664
rect 45373 56661 45385 56664
rect 45419 56661 45431 56695
rect 48222 56692 48228 56704
rect 48183 56664 48228 56692
rect 45373 56655 45431 56661
rect 48222 56652 48228 56664
rect 48280 56652 48286 56704
rect 50154 56692 50160 56704
rect 50115 56664 50160 56692
rect 50154 56652 50160 56664
rect 50212 56652 50218 56704
rect 67082 56652 67088 56704
rect 67140 56692 67146 56704
rect 67284 56701 67312 56732
rect 67913 56729 67925 56732
rect 67959 56729 67971 56763
rect 67913 56723 67971 56729
rect 67269 56695 67327 56701
rect 67269 56692 67281 56695
rect 67140 56664 67281 56692
rect 67140 56652 67146 56664
rect 67269 56661 67281 56664
rect 67315 56661 67327 56695
rect 67269 56655 67327 56661
rect 1104 56602 68816 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 68816 56602
rect 1104 56528 68816 56550
rect 2130 56448 2136 56500
rect 2188 56488 2194 56500
rect 26142 56488 26148 56500
rect 2188 56460 26004 56488
rect 26103 56460 26148 56488
rect 2188 56448 2194 56460
rect 16942 56429 16948 56432
rect 16936 56420 16948 56429
rect 16903 56392 16948 56420
rect 16936 56383 16948 56392
rect 16942 56380 16948 56383
rect 17000 56380 17006 56432
rect 19972 56423 20030 56429
rect 19972 56389 19984 56423
rect 20018 56420 20030 56423
rect 20346 56420 20352 56432
rect 20018 56392 20352 56420
rect 20018 56389 20030 56392
rect 19972 56383 20030 56389
rect 20346 56380 20352 56392
rect 20404 56380 20410 56432
rect 25976 56420 26004 56460
rect 26142 56448 26148 56460
rect 26200 56448 26206 56500
rect 28534 56448 28540 56500
rect 28592 56488 28598 56500
rect 29638 56488 29644 56500
rect 28592 56460 29644 56488
rect 28592 56448 28598 56460
rect 29638 56448 29644 56460
rect 29696 56448 29702 56500
rect 30837 56491 30895 56497
rect 30837 56457 30849 56491
rect 30883 56488 30895 56491
rect 30926 56488 30932 56500
rect 30883 56460 30932 56488
rect 30883 56457 30895 56460
rect 30837 56451 30895 56457
rect 30926 56448 30932 56460
rect 30984 56448 30990 56500
rect 35066 56448 35072 56500
rect 35124 56488 35130 56500
rect 35805 56491 35863 56497
rect 35805 56488 35817 56491
rect 35124 56460 35817 56488
rect 35124 56448 35130 56460
rect 35805 56457 35817 56460
rect 35851 56457 35863 56491
rect 35805 56451 35863 56457
rect 37366 56448 37372 56500
rect 37424 56488 37430 56500
rect 40678 56488 40684 56500
rect 37424 56460 40684 56488
rect 37424 56448 37430 56460
rect 40678 56448 40684 56460
rect 40736 56448 40742 56500
rect 40865 56491 40923 56497
rect 40865 56457 40877 56491
rect 40911 56488 40923 56491
rect 41322 56488 41328 56500
rect 40911 56460 41328 56488
rect 40911 56457 40923 56460
rect 40865 56451 40923 56457
rect 41322 56448 41328 56460
rect 41380 56448 41386 56500
rect 43346 56488 43352 56500
rect 43307 56460 43352 56488
rect 43346 56448 43352 56460
rect 43404 56448 43410 56500
rect 26878 56420 26884 56432
rect 25976 56392 26884 56420
rect 26878 56380 26884 56392
rect 26936 56380 26942 56432
rect 27522 56380 27528 56432
rect 27580 56420 27586 56432
rect 27580 56392 28672 56420
rect 27580 56380 27586 56392
rect 15105 56355 15163 56361
rect 15105 56321 15117 56355
rect 15151 56352 15163 56355
rect 15378 56352 15384 56364
rect 15151 56324 15384 56352
rect 15151 56321 15163 56324
rect 15105 56315 15163 56321
rect 15378 56312 15384 56324
rect 15436 56312 15442 56364
rect 19426 56312 19432 56364
rect 19484 56352 19490 56364
rect 19705 56355 19763 56361
rect 19705 56352 19717 56355
rect 19484 56324 19717 56352
rect 19484 56312 19490 56324
rect 19705 56321 19717 56324
rect 19751 56321 19763 56355
rect 19705 56315 19763 56321
rect 21726 56312 21732 56364
rect 21784 56352 21790 56364
rect 22005 56355 22063 56361
rect 22005 56352 22017 56355
rect 21784 56324 22017 56352
rect 21784 56312 21790 56324
rect 22005 56321 22017 56324
rect 22051 56321 22063 56355
rect 22186 56352 22192 56364
rect 22147 56324 22192 56352
rect 22005 56315 22063 56321
rect 22186 56312 22192 56324
rect 22244 56312 22250 56364
rect 22281 56355 22339 56361
rect 22281 56321 22293 56355
rect 22327 56352 22339 56355
rect 22370 56352 22376 56364
rect 22327 56324 22376 56352
rect 22327 56321 22339 56324
rect 22281 56315 22339 56321
rect 22370 56312 22376 56324
rect 22428 56312 22434 56364
rect 24765 56355 24823 56361
rect 24765 56321 24777 56355
rect 24811 56352 24823 56355
rect 24946 56352 24952 56364
rect 24811 56324 24952 56352
rect 24811 56321 24823 56324
rect 24765 56315 24823 56321
rect 24946 56312 24952 56324
rect 25004 56312 25010 56364
rect 25406 56312 25412 56364
rect 25464 56352 25470 56364
rect 25501 56355 25559 56361
rect 25501 56352 25513 56355
rect 25464 56324 25513 56352
rect 25464 56312 25470 56324
rect 25501 56321 25513 56324
rect 25547 56321 25559 56355
rect 25501 56315 25559 56321
rect 26145 56355 26203 56361
rect 26145 56321 26157 56355
rect 26191 56352 26203 56355
rect 26418 56352 26424 56364
rect 26191 56324 26424 56352
rect 26191 56321 26203 56324
rect 26145 56315 26203 56321
rect 26418 56312 26424 56324
rect 26476 56312 26482 56364
rect 27424 56355 27482 56361
rect 27424 56321 27436 56355
rect 27470 56352 27482 56355
rect 28534 56352 28540 56364
rect 27470 56324 28540 56352
rect 27470 56321 27482 56324
rect 27424 56315 27482 56321
rect 28534 56312 28540 56324
rect 28592 56312 28598 56364
rect 28644 56352 28672 56392
rect 33318 56380 33324 56432
rect 33376 56420 33382 56432
rect 33566 56423 33624 56429
rect 33566 56420 33578 56423
rect 33376 56392 33578 56420
rect 33376 56380 33382 56392
rect 33566 56389 33578 56392
rect 33612 56389 33624 56423
rect 33566 56383 33624 56389
rect 35437 56423 35495 56429
rect 35437 56389 35449 56423
rect 35483 56420 35495 56423
rect 36722 56420 36728 56432
rect 35483 56392 36728 56420
rect 35483 56389 35495 56392
rect 35437 56383 35495 56389
rect 36722 56380 36728 56392
rect 36780 56380 36786 56432
rect 42886 56420 42892 56432
rect 42628 56392 42892 56420
rect 35529 56355 35587 56361
rect 28644 56324 29316 56352
rect 16022 56244 16028 56296
rect 16080 56284 16086 56296
rect 16669 56287 16727 56293
rect 16669 56284 16681 56287
rect 16080 56256 16681 56284
rect 16080 56244 16086 56256
rect 16669 56253 16681 56256
rect 16715 56253 16727 56287
rect 27154 56284 27160 56296
rect 27115 56256 27160 56284
rect 16669 56247 16727 56253
rect 27154 56244 27160 56256
rect 27212 56244 27218 56296
rect 28997 56287 29055 56293
rect 28997 56284 29009 56287
rect 28552 56256 29009 56284
rect 14918 56216 14924 56228
rect 14879 56188 14924 56216
rect 14918 56176 14924 56188
rect 14976 56176 14982 56228
rect 18049 56219 18107 56225
rect 18049 56185 18061 56219
rect 18095 56216 18107 56219
rect 18138 56216 18144 56228
rect 18095 56188 18144 56216
rect 18095 56185 18107 56188
rect 18049 56179 18107 56185
rect 18138 56176 18144 56188
rect 18196 56176 18202 56228
rect 28442 56176 28448 56228
rect 28500 56216 28506 56228
rect 28552 56225 28580 56256
rect 28997 56253 29009 56256
rect 29043 56253 29055 56287
rect 29181 56287 29239 56293
rect 29181 56284 29193 56287
rect 28997 56247 29055 56253
rect 29104 56256 29193 56284
rect 28537 56219 28595 56225
rect 28537 56216 28549 56219
rect 28500 56188 28549 56216
rect 28500 56176 28506 56188
rect 28537 56185 28549 56188
rect 28583 56185 28595 56219
rect 28537 56179 28595 56185
rect 19334 56108 19340 56160
rect 19392 56148 19398 56160
rect 21085 56151 21143 56157
rect 21085 56148 21097 56151
rect 19392 56120 21097 56148
rect 19392 56108 19398 56120
rect 21085 56117 21097 56120
rect 21131 56117 21143 56151
rect 21085 56111 21143 56117
rect 21821 56151 21879 56157
rect 21821 56117 21833 56151
rect 21867 56148 21879 56151
rect 22738 56148 22744 56160
rect 21867 56120 22744 56148
rect 21867 56117 21879 56120
rect 21821 56111 21879 56117
rect 22738 56108 22744 56120
rect 22796 56108 22802 56160
rect 24486 56108 24492 56160
rect 24544 56148 24550 56160
rect 24581 56151 24639 56157
rect 24581 56148 24593 56151
rect 24544 56120 24593 56148
rect 24544 56108 24550 56120
rect 24581 56117 24593 56120
rect 24627 56117 24639 56151
rect 25314 56148 25320 56160
rect 25275 56120 25320 56148
rect 24581 56111 24639 56117
rect 25314 56108 25320 56120
rect 25372 56108 25378 56160
rect 29104 56148 29132 56256
rect 29181 56253 29193 56256
rect 29227 56253 29239 56287
rect 29288 56284 29316 56324
rect 35529 56321 35541 56355
rect 35575 56321 35587 56355
rect 35529 56315 35587 56321
rect 35621 56355 35679 56361
rect 35621 56321 35633 56355
rect 35667 56352 35679 56355
rect 36170 56352 36176 56364
rect 35667 56324 36176 56352
rect 35667 56321 35679 56324
rect 35621 56315 35679 56321
rect 30098 56293 30104 56296
rect 29917 56287 29975 56293
rect 29917 56284 29929 56287
rect 29288 56256 29929 56284
rect 29181 56247 29239 56253
rect 29917 56253 29929 56256
rect 29963 56253 29975 56287
rect 29917 56247 29975 56253
rect 30055 56287 30104 56293
rect 30055 56253 30067 56287
rect 30101 56253 30104 56287
rect 30055 56247 30104 56253
rect 30098 56244 30104 56247
rect 30156 56244 30162 56296
rect 30190 56244 30196 56296
rect 30248 56284 30254 56296
rect 30248 56256 30293 56284
rect 30248 56244 30254 56256
rect 33042 56244 33048 56296
rect 33100 56284 33106 56296
rect 33321 56287 33379 56293
rect 33321 56284 33333 56287
rect 33100 56256 33333 56284
rect 33100 56244 33106 56256
rect 33321 56253 33333 56256
rect 33367 56253 33379 56287
rect 35544 56284 35572 56315
rect 36170 56312 36176 56324
rect 36228 56312 36234 56364
rect 36357 56355 36415 56361
rect 36357 56321 36369 56355
rect 36403 56352 36415 56355
rect 37366 56352 37372 56364
rect 36403 56324 37372 56352
rect 36403 56321 36415 56324
rect 36357 56315 36415 56321
rect 37366 56312 37372 56324
rect 37424 56312 37430 56364
rect 38746 56312 38752 56364
rect 38804 56352 38810 56364
rect 39209 56355 39267 56361
rect 39209 56352 39221 56355
rect 38804 56324 39221 56352
rect 38804 56312 38810 56324
rect 39209 56321 39221 56324
rect 39255 56321 39267 56355
rect 39209 56315 39267 56321
rect 39301 56355 39359 56361
rect 39301 56321 39313 56355
rect 39347 56321 39359 56355
rect 39301 56315 39359 56321
rect 39393 56355 39451 56361
rect 39393 56321 39405 56355
rect 39439 56321 39451 56355
rect 40494 56352 40500 56364
rect 40455 56324 40500 56352
rect 39393 56315 39451 56321
rect 35986 56284 35992 56296
rect 35544 56256 35992 56284
rect 33321 56247 33379 56253
rect 35986 56244 35992 56256
rect 36044 56244 36050 56296
rect 36188 56284 36216 56312
rect 37182 56284 37188 56296
rect 36188 56256 37188 56284
rect 37182 56244 37188 56256
rect 37240 56284 37246 56296
rect 38838 56284 38844 56296
rect 37240 56256 38844 56284
rect 37240 56244 37246 56256
rect 38838 56244 38844 56256
rect 38896 56284 38902 56296
rect 39316 56284 39344 56315
rect 38896 56256 39344 56284
rect 39408 56284 39436 56315
rect 40494 56312 40500 56324
rect 40552 56312 40558 56364
rect 40678 56352 40684 56364
rect 40639 56324 40684 56352
rect 40678 56312 40684 56324
rect 40736 56312 40742 56364
rect 42628 56361 42656 56392
rect 42886 56380 42892 56392
rect 42944 56380 42950 56432
rect 49412 56423 49470 56429
rect 49412 56389 49424 56423
rect 49458 56420 49470 56423
rect 50154 56420 50160 56432
rect 49458 56392 50160 56420
rect 49458 56389 49470 56392
rect 49412 56383 49470 56389
rect 50154 56380 50160 56392
rect 50212 56380 50218 56432
rect 42613 56355 42671 56361
rect 42613 56321 42625 56355
rect 42659 56321 42671 56355
rect 43530 56352 43536 56364
rect 43491 56324 43536 56352
rect 42613 56315 42671 56321
rect 43530 56312 43536 56324
rect 43588 56312 43594 56364
rect 45186 56352 45192 56364
rect 45147 56324 45192 56352
rect 45186 56312 45192 56324
rect 45244 56312 45250 56364
rect 45456 56355 45514 56361
rect 45456 56321 45468 56355
rect 45502 56352 45514 56355
rect 45830 56352 45836 56364
rect 45502 56324 45836 56352
rect 45502 56321 45514 56324
rect 45456 56315 45514 56321
rect 45830 56312 45836 56324
rect 45888 56312 45894 56364
rect 48222 56352 48228 56364
rect 48183 56324 48228 56352
rect 48222 56312 48228 56324
rect 48280 56312 48286 56364
rect 48317 56355 48375 56361
rect 48317 56321 48329 56355
rect 48363 56352 48375 56355
rect 49694 56352 49700 56364
rect 48363 56324 49700 56352
rect 48363 56321 48375 56324
rect 48317 56315 48375 56321
rect 49694 56312 49700 56324
rect 49752 56352 49758 56364
rect 50338 56352 50344 56364
rect 49752 56324 50344 56352
rect 49752 56312 49758 56324
rect 50338 56312 50344 56324
rect 50396 56312 50402 56364
rect 39408 56256 42104 56284
rect 38896 56244 38902 56256
rect 29638 56216 29644 56228
rect 29599 56188 29644 56216
rect 29638 56176 29644 56188
rect 29696 56176 29702 56228
rect 34606 56176 34612 56228
rect 34664 56216 34670 56228
rect 35253 56219 35311 56225
rect 35253 56216 35265 56219
rect 34664 56188 35265 56216
rect 34664 56176 34670 56188
rect 35253 56185 35265 56188
rect 35299 56185 35311 56219
rect 36004 56216 36032 56244
rect 36630 56216 36636 56228
rect 36004 56188 36636 56216
rect 35253 56179 35311 56185
rect 36630 56176 36636 56188
rect 36688 56176 36694 56228
rect 38194 56176 38200 56228
rect 38252 56216 38258 56228
rect 39025 56219 39083 56225
rect 39025 56216 39037 56219
rect 38252 56188 39037 56216
rect 38252 56176 38258 56188
rect 39025 56185 39037 56188
rect 39071 56185 39083 56219
rect 39025 56179 39083 56185
rect 39577 56219 39635 56225
rect 39577 56185 39589 56219
rect 39623 56216 39635 56219
rect 41598 56216 41604 56228
rect 39623 56188 41604 56216
rect 39623 56185 39635 56188
rect 39577 56179 39635 56185
rect 41598 56176 41604 56188
rect 41656 56176 41662 56228
rect 42076 56216 42104 56256
rect 42150 56244 42156 56296
rect 42208 56284 42214 56296
rect 42794 56284 42800 56296
rect 42208 56256 42800 56284
rect 42208 56244 42214 56256
rect 42794 56244 42800 56256
rect 42852 56284 42858 56296
rect 42889 56287 42947 56293
rect 42889 56284 42901 56287
rect 42852 56256 42901 56284
rect 42852 56244 42858 56256
rect 42889 56253 42901 56256
rect 42935 56253 42947 56287
rect 42889 56247 42947 56253
rect 43809 56287 43867 56293
rect 43809 56253 43821 56287
rect 43855 56284 43867 56287
rect 43898 56284 43904 56296
rect 43855 56256 43904 56284
rect 43855 56253 43867 56256
rect 43809 56247 43867 56253
rect 43898 56244 43904 56256
rect 43956 56244 43962 56296
rect 48774 56244 48780 56296
rect 48832 56284 48838 56296
rect 49145 56287 49203 56293
rect 49145 56284 49157 56287
rect 48832 56256 49157 56284
rect 48832 56244 48838 56256
rect 49145 56253 49157 56256
rect 49191 56253 49203 56287
rect 49145 56247 49203 56253
rect 42610 56216 42616 56228
rect 42076 56188 42616 56216
rect 42610 56176 42616 56188
rect 42668 56216 42674 56228
rect 43717 56219 43775 56225
rect 43717 56216 43729 56219
rect 42668 56188 43729 56216
rect 42668 56176 42674 56188
rect 43717 56185 43729 56188
rect 43763 56185 43775 56219
rect 43717 56179 43775 56185
rect 30374 56148 30380 56160
rect 29104 56120 30380 56148
rect 30374 56108 30380 56120
rect 30432 56108 30438 56160
rect 32306 56108 32312 56160
rect 32364 56148 32370 56160
rect 34701 56151 34759 56157
rect 34701 56148 34713 56151
rect 32364 56120 34713 56148
rect 32364 56108 32370 56120
rect 34701 56117 34713 56120
rect 34747 56148 34759 56151
rect 35802 56148 35808 56160
rect 34747 56120 35808 56148
rect 34747 56117 34759 56120
rect 34701 56111 34759 56117
rect 35802 56108 35808 56120
rect 35860 56108 35866 56160
rect 35894 56108 35900 56160
rect 35952 56148 35958 56160
rect 36541 56151 36599 56157
rect 36541 56148 36553 56151
rect 35952 56120 36553 56148
rect 35952 56108 35958 56120
rect 36541 56117 36553 56120
rect 36587 56148 36599 56151
rect 37090 56148 37096 56160
rect 36587 56120 37096 56148
rect 36587 56117 36599 56120
rect 36541 56111 36599 56117
rect 37090 56108 37096 56120
rect 37148 56108 37154 56160
rect 42426 56148 42432 56160
rect 42387 56120 42432 56148
rect 42426 56108 42432 56120
rect 42484 56108 42490 56160
rect 42797 56151 42855 56157
rect 42797 56117 42809 56151
rect 42843 56148 42855 56151
rect 42978 56148 42984 56160
rect 42843 56120 42984 56148
rect 42843 56117 42855 56120
rect 42797 56111 42855 56117
rect 42978 56108 42984 56120
rect 43036 56108 43042 56160
rect 46566 56148 46572 56160
rect 46527 56120 46572 56148
rect 46566 56108 46572 56120
rect 46624 56108 46630 56160
rect 47762 56108 47768 56160
rect 47820 56148 47826 56160
rect 48501 56151 48559 56157
rect 48501 56148 48513 56151
rect 47820 56120 48513 56148
rect 47820 56108 47826 56120
rect 48501 56117 48513 56120
rect 48547 56117 48559 56151
rect 50522 56148 50528 56160
rect 50483 56120 50528 56148
rect 48501 56111 48559 56117
rect 50522 56108 50528 56120
rect 50580 56108 50586 56160
rect 1104 56058 68816 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 65654 56058
rect 65706 56006 65718 56058
rect 65770 56006 65782 56058
rect 65834 56006 65846 56058
rect 65898 56006 65910 56058
rect 65962 56006 68816 56058
rect 1104 55984 68816 56006
rect 16022 55944 16028 55956
rect 15983 55916 16028 55944
rect 16022 55904 16028 55916
rect 16080 55904 16086 55956
rect 20073 55947 20131 55953
rect 20073 55913 20085 55947
rect 20119 55913 20131 55947
rect 20073 55907 20131 55913
rect 20257 55947 20315 55953
rect 20257 55913 20269 55947
rect 20303 55944 20315 55947
rect 20530 55944 20536 55956
rect 20303 55916 20536 55944
rect 20303 55913 20315 55916
rect 20257 55907 20315 55913
rect 20088 55876 20116 55907
rect 20530 55904 20536 55916
rect 20588 55904 20594 55956
rect 22830 55904 22836 55956
rect 22888 55944 22894 55956
rect 23201 55947 23259 55953
rect 23201 55944 23213 55947
rect 22888 55916 23213 55944
rect 22888 55904 22894 55916
rect 23201 55913 23213 55916
rect 23247 55913 23259 55947
rect 26510 55944 26516 55956
rect 26471 55916 26516 55944
rect 23201 55907 23259 55913
rect 26510 55904 26516 55916
rect 26568 55904 26574 55956
rect 26878 55904 26884 55956
rect 26936 55944 26942 55956
rect 26936 55916 30144 55944
rect 26936 55904 26942 55916
rect 20438 55876 20444 55888
rect 20088 55848 20444 55876
rect 20438 55836 20444 55848
rect 20496 55836 20502 55888
rect 29917 55879 29975 55885
rect 29917 55845 29929 55879
rect 29963 55876 29975 55879
rect 30006 55876 30012 55888
rect 29963 55848 30012 55876
rect 29963 55845 29975 55848
rect 29917 55839 29975 55845
rect 30006 55836 30012 55848
rect 30064 55836 30070 55888
rect 30116 55876 30144 55916
rect 30282 55904 30288 55956
rect 30340 55944 30346 55956
rect 30561 55947 30619 55953
rect 30561 55944 30573 55947
rect 30340 55916 30573 55944
rect 30340 55904 30346 55916
rect 30561 55913 30573 55916
rect 30607 55913 30619 55947
rect 30561 55907 30619 55913
rect 30834 55904 30840 55956
rect 30892 55944 30898 55956
rect 31205 55947 31263 55953
rect 31205 55944 31217 55947
rect 30892 55916 31217 55944
rect 30892 55904 30898 55916
rect 31205 55913 31217 55916
rect 31251 55913 31263 55947
rect 36814 55944 36820 55956
rect 31205 55907 31263 55913
rect 35820 55916 36820 55944
rect 34606 55876 34612 55888
rect 30116 55848 34612 55876
rect 34606 55836 34612 55848
rect 34664 55876 34670 55888
rect 34664 55848 35112 55876
rect 34664 55836 34670 55848
rect 24486 55808 24492 55820
rect 24447 55780 24492 55808
rect 24486 55768 24492 55780
rect 24544 55768 24550 55820
rect 27525 55811 27583 55817
rect 27525 55808 27537 55811
rect 26712 55780 27537 55808
rect 14829 55743 14887 55749
rect 14829 55709 14841 55743
rect 14875 55740 14887 55743
rect 15286 55740 15292 55752
rect 14875 55712 15292 55740
rect 14875 55709 14887 55712
rect 14829 55703 14887 55709
rect 15286 55700 15292 55712
rect 15344 55700 15350 55752
rect 16025 55743 16083 55749
rect 16025 55709 16037 55743
rect 16071 55740 16083 55743
rect 16761 55743 16819 55749
rect 16761 55740 16773 55743
rect 16071 55712 16773 55740
rect 16071 55709 16083 55712
rect 16025 55703 16083 55709
rect 16761 55709 16773 55712
rect 16807 55740 16819 55743
rect 17310 55740 17316 55752
rect 16807 55712 17316 55740
rect 16807 55709 16819 55712
rect 16761 55703 16819 55709
rect 17310 55700 17316 55712
rect 17368 55700 17374 55752
rect 21821 55743 21879 55749
rect 21821 55709 21833 55743
rect 21867 55740 21879 55743
rect 23198 55740 23204 55752
rect 21867 55712 23204 55740
rect 21867 55709 21879 55712
rect 21821 55703 21879 55709
rect 23198 55700 23204 55712
rect 23256 55700 23262 55752
rect 24756 55743 24814 55749
rect 24756 55709 24768 55743
rect 24802 55740 24814 55743
rect 25314 55740 25320 55752
rect 24802 55712 25320 55740
rect 24802 55709 24814 55712
rect 24756 55703 24814 55709
rect 25314 55700 25320 55712
rect 25372 55700 25378 55752
rect 26712 55749 26740 55780
rect 27525 55777 27537 55780
rect 27571 55777 27583 55811
rect 28442 55808 28448 55820
rect 28403 55780 28448 55808
rect 27525 55771 27583 55777
rect 28442 55768 28448 55780
rect 28500 55768 28506 55820
rect 34790 55808 34796 55820
rect 29748 55780 34796 55808
rect 26697 55743 26755 55749
rect 26697 55709 26709 55743
rect 26743 55709 26755 55743
rect 26697 55703 26755 55709
rect 27249 55743 27307 55749
rect 27249 55709 27261 55743
rect 27295 55709 27307 55743
rect 27249 55703 27307 55709
rect 27341 55743 27399 55749
rect 27341 55709 27353 55743
rect 27387 55740 27399 55743
rect 27614 55740 27620 55752
rect 27387 55712 27620 55740
rect 27387 55709 27399 55712
rect 27341 55703 27399 55709
rect 19334 55632 19340 55684
rect 19392 55672 19398 55684
rect 19889 55675 19947 55681
rect 19889 55672 19901 55675
rect 19392 55644 19901 55672
rect 19392 55632 19398 55644
rect 19889 55641 19901 55644
rect 19935 55641 19947 55675
rect 19889 55635 19947 55641
rect 22088 55675 22146 55681
rect 22088 55641 22100 55675
rect 22134 55672 22146 55675
rect 22186 55672 22192 55684
rect 22134 55644 22192 55672
rect 22134 55641 22146 55644
rect 22088 55635 22146 55641
rect 22186 55632 22192 55644
rect 22244 55632 22250 55684
rect 27264 55672 27292 55703
rect 27614 55700 27620 55712
rect 27672 55700 27678 55752
rect 28350 55700 28356 55752
rect 28408 55740 28414 55752
rect 29748 55749 29776 55780
rect 34790 55768 34796 55780
rect 34848 55768 34854 55820
rect 28629 55743 28687 55749
rect 28629 55740 28641 55743
rect 28408 55712 28641 55740
rect 28408 55700 28414 55712
rect 28629 55709 28641 55712
rect 28675 55709 28687 55743
rect 28629 55703 28687 55709
rect 29733 55743 29791 55749
rect 29733 55709 29745 55743
rect 29779 55709 29791 55743
rect 29733 55703 29791 55709
rect 29822 55700 29828 55752
rect 29880 55740 29886 55752
rect 30558 55740 30564 55752
rect 29880 55712 30564 55740
rect 29880 55700 29886 55712
rect 30558 55700 30564 55712
rect 30616 55740 30622 55752
rect 31205 55743 31263 55749
rect 31205 55740 31217 55743
rect 30616 55712 31217 55740
rect 30616 55700 30622 55712
rect 31205 55709 31217 55712
rect 31251 55709 31263 55743
rect 32306 55740 32312 55752
rect 32267 55712 32312 55740
rect 31205 55703 31263 55709
rect 32306 55700 32312 55712
rect 32364 55700 32370 55752
rect 35084 55740 35112 55848
rect 35820 55740 35848 55916
rect 36814 55904 36820 55916
rect 36872 55904 36878 55956
rect 45830 55944 45836 55956
rect 36924 55916 43484 55944
rect 45791 55916 45836 55944
rect 36924 55885 36952 55916
rect 36909 55879 36967 55885
rect 36909 55876 36921 55879
rect 36004 55848 36921 55876
rect 36004 55749 36032 55848
rect 36909 55845 36921 55848
rect 36955 55845 36967 55879
rect 36909 55839 36967 55845
rect 38197 55879 38255 55885
rect 38197 55845 38209 55879
rect 38243 55876 38255 55879
rect 43456 55876 43484 55916
rect 45830 55904 45836 55916
rect 45888 55904 45894 55956
rect 46842 55944 46848 55956
rect 46803 55916 46848 55944
rect 46842 55904 46848 55916
rect 46900 55904 46906 55956
rect 46934 55904 46940 55956
rect 46992 55944 46998 55956
rect 48590 55944 48596 55956
rect 46992 55916 48596 55944
rect 46992 55904 46998 55916
rect 48590 55904 48596 55916
rect 48648 55904 48654 55956
rect 48774 55944 48780 55956
rect 48735 55916 48780 55944
rect 48774 55904 48780 55916
rect 48832 55904 48838 55956
rect 50525 55947 50583 55953
rect 50525 55913 50537 55947
rect 50571 55944 50583 55947
rect 50614 55944 50620 55956
rect 50571 55916 50620 55944
rect 50571 55913 50583 55916
rect 50525 55907 50583 55913
rect 50614 55904 50620 55916
rect 50672 55904 50678 55956
rect 55674 55876 55680 55888
rect 38243 55848 38884 55876
rect 43456 55848 46704 55876
rect 38243 55845 38255 55848
rect 38197 55839 38255 55845
rect 36078 55768 36084 55820
rect 36136 55808 36142 55820
rect 36449 55811 36507 55817
rect 36449 55808 36461 55811
rect 36136 55780 36461 55808
rect 36136 55768 36142 55780
rect 36449 55777 36461 55780
rect 36495 55777 36507 55811
rect 36449 55771 36507 55777
rect 36630 55768 36636 55820
rect 36688 55808 36694 55820
rect 38746 55808 38752 55820
rect 36688 55780 38752 55808
rect 36688 55768 36694 55780
rect 35084 55712 35848 55740
rect 27522 55672 27528 55684
rect 27264 55644 27528 55672
rect 27522 55632 27528 55644
rect 27580 55632 27586 55684
rect 30098 55672 30104 55684
rect 27632 55644 30104 55672
rect 14642 55604 14648 55616
rect 14603 55576 14648 55604
rect 14642 55564 14648 55576
rect 14700 55564 14706 55616
rect 16761 55607 16819 55613
rect 16761 55573 16773 55607
rect 16807 55604 16819 55607
rect 16942 55604 16948 55616
rect 16807 55576 16948 55604
rect 16807 55573 16819 55576
rect 16761 55567 16819 55573
rect 16942 55564 16948 55576
rect 17000 55564 17006 55616
rect 20070 55564 20076 55616
rect 20128 55613 20134 55616
rect 20128 55607 20147 55613
rect 20135 55573 20147 55607
rect 20128 55567 20147 55573
rect 20128 55564 20134 55567
rect 25130 55564 25136 55616
rect 25188 55604 25194 55616
rect 25869 55607 25927 55613
rect 25869 55604 25881 55607
rect 25188 55576 25881 55604
rect 25188 55564 25194 55576
rect 25869 55573 25881 55576
rect 25915 55604 25927 55607
rect 27632 55604 27660 55644
rect 30098 55632 30104 55644
rect 30156 55632 30162 55684
rect 30374 55672 30380 55684
rect 30335 55644 30380 55672
rect 30374 55632 30380 55644
rect 30432 55632 30438 55684
rect 32493 55675 32551 55681
rect 32493 55641 32505 55675
rect 32539 55672 32551 55675
rect 32674 55672 32680 55684
rect 32539 55644 32680 55672
rect 32539 55641 32551 55644
rect 32493 55635 32551 55641
rect 32674 55632 32680 55644
rect 32732 55632 32738 55684
rect 34146 55672 34152 55684
rect 34107 55644 34152 55672
rect 34146 55632 34152 55644
rect 34204 55632 34210 55684
rect 25915 55576 27660 55604
rect 25915 55573 25927 55576
rect 25869 55567 25927 55573
rect 28718 55564 28724 55616
rect 28776 55604 28782 55616
rect 28813 55607 28871 55613
rect 28813 55604 28825 55607
rect 28776 55576 28825 55604
rect 28776 55564 28782 55576
rect 28813 55573 28825 55576
rect 28859 55573 28871 55607
rect 28813 55567 28871 55573
rect 29730 55564 29736 55616
rect 29788 55604 29794 55616
rect 30466 55604 30472 55616
rect 29788 55576 30472 55604
rect 29788 55564 29794 55576
rect 30466 55564 30472 55576
rect 30524 55604 30530 55616
rect 30577 55607 30635 55613
rect 30577 55604 30589 55607
rect 30524 55576 30589 55604
rect 30524 55564 30530 55576
rect 30577 55573 30589 55576
rect 30623 55573 30635 55607
rect 30742 55604 30748 55616
rect 30703 55576 30748 55604
rect 30577 55567 30635 55573
rect 30742 55564 30748 55576
rect 30800 55564 30806 55616
rect 34606 55564 34612 55616
rect 34664 55604 34670 55616
rect 35713 55607 35771 55613
rect 35713 55604 35725 55607
rect 34664 55576 35725 55604
rect 34664 55564 34670 55576
rect 35713 55573 35725 55576
rect 35759 55573 35771 55607
rect 35820 55604 35848 55712
rect 35989 55743 36047 55749
rect 35989 55709 36001 55743
rect 36035 55709 36047 55743
rect 35989 55703 36047 55709
rect 36262 55700 36268 55752
rect 36320 55740 36326 55752
rect 36357 55743 36415 55749
rect 36357 55740 36369 55743
rect 36320 55712 36369 55740
rect 36320 55700 36326 55712
rect 36357 55709 36369 55712
rect 36403 55709 36415 55743
rect 36357 55703 36415 55709
rect 36814 55700 36820 55752
rect 36872 55740 36878 55752
rect 37093 55743 37151 55749
rect 37093 55740 37105 55743
rect 36872 55712 37105 55740
rect 36872 55700 36878 55712
rect 37093 55709 37105 55712
rect 37139 55709 37151 55743
rect 37093 55703 37151 55709
rect 37182 55700 37188 55752
rect 37240 55740 37246 55752
rect 37461 55743 37519 55749
rect 37240 55712 37412 55740
rect 37240 55700 37246 55712
rect 35894 55632 35900 55684
rect 35952 55672 35958 55684
rect 37277 55675 37335 55681
rect 37277 55672 37289 55675
rect 35952 55644 37289 55672
rect 35952 55632 35958 55644
rect 37277 55641 37289 55644
rect 37323 55641 37335 55675
rect 37384 55672 37412 55712
rect 37461 55709 37473 55743
rect 37507 55740 37519 55743
rect 38194 55740 38200 55752
rect 37507 55712 38200 55740
rect 37507 55709 37519 55712
rect 37461 55703 37519 55709
rect 38194 55700 38200 55712
rect 38252 55700 38258 55752
rect 37921 55675 37979 55681
rect 37921 55672 37933 55675
rect 37384 55644 37933 55672
rect 37277 55635 37335 55641
rect 37921 55641 37933 55644
rect 37967 55641 37979 55675
rect 37921 55635 37979 55641
rect 38105 55675 38163 55681
rect 38105 55641 38117 55675
rect 38151 55672 38163 55675
rect 38304 55672 38332 55780
rect 38746 55768 38752 55780
rect 38804 55768 38810 55820
rect 38856 55817 38884 55848
rect 38841 55811 38899 55817
rect 38841 55777 38853 55811
rect 38887 55808 38899 55811
rect 39114 55808 39120 55820
rect 38887 55780 39120 55808
rect 38887 55777 38899 55780
rect 38841 55771 38899 55777
rect 39114 55768 39120 55780
rect 39172 55768 39178 55820
rect 45005 55811 45063 55817
rect 45005 55777 45017 55811
rect 45051 55808 45063 55811
rect 46566 55808 46572 55820
rect 45051 55780 46572 55808
rect 45051 55777 45063 55780
rect 45005 55771 45063 55777
rect 46566 55768 46572 55780
rect 46624 55768 46630 55820
rect 46676 55808 46704 55848
rect 47320 55848 55680 55876
rect 47320 55808 47348 55848
rect 55674 55836 55680 55848
rect 55732 55836 55738 55888
rect 46676 55780 47348 55808
rect 47673 55811 47731 55817
rect 47673 55777 47685 55811
rect 47719 55808 47731 55811
rect 48222 55808 48228 55820
rect 47719 55780 48228 55808
rect 47719 55777 47731 55780
rect 47673 55771 47731 55777
rect 48222 55768 48228 55780
rect 48280 55768 48286 55820
rect 50157 55811 50215 55817
rect 50157 55808 50169 55811
rect 48516 55780 50169 55808
rect 38930 55740 38936 55752
rect 38891 55712 38936 55740
rect 38930 55700 38936 55712
rect 38988 55700 38994 55752
rect 39022 55700 39028 55752
rect 39080 55740 39086 55752
rect 40129 55743 40187 55749
rect 39080 55712 39620 55740
rect 39080 55700 39086 55712
rect 38151 55644 38332 55672
rect 38151 55641 38163 55644
rect 38105 55635 38163 55641
rect 36081 55607 36139 55613
rect 36081 55604 36093 55607
rect 35820 55576 36093 55604
rect 35713 55567 35771 55573
rect 36081 55573 36093 55576
rect 36127 55573 36139 55607
rect 36081 55567 36139 55573
rect 36173 55607 36231 55613
rect 36173 55573 36185 55607
rect 36219 55604 36231 55607
rect 36630 55604 36636 55616
rect 36219 55576 36636 55604
rect 36219 55573 36231 55576
rect 36173 55567 36231 55573
rect 36630 55564 36636 55576
rect 36688 55564 36694 55616
rect 37182 55604 37188 55616
rect 37143 55576 37188 55604
rect 37182 55564 37188 55576
rect 37240 55564 37246 55616
rect 38654 55604 38660 55616
rect 38615 55576 38660 55604
rect 38654 55564 38660 55576
rect 38712 55564 38718 55616
rect 39592 55604 39620 55712
rect 40129 55709 40141 55743
rect 40175 55740 40187 55743
rect 40770 55740 40776 55752
rect 40175 55712 40776 55740
rect 40175 55709 40187 55712
rect 40129 55703 40187 55709
rect 40770 55700 40776 55712
rect 40828 55700 40834 55752
rect 45186 55740 45192 55752
rect 45147 55712 45192 55740
rect 45186 55700 45192 55712
rect 45244 55700 45250 55752
rect 45373 55743 45431 55749
rect 45373 55709 45385 55743
rect 45419 55740 45431 55743
rect 46017 55743 46075 55749
rect 46017 55740 46029 55743
rect 45419 55712 46029 55740
rect 45419 55709 45431 55712
rect 45373 55703 45431 55709
rect 46017 55709 46029 55712
rect 46063 55709 46075 55743
rect 46017 55703 46075 55709
rect 40396 55675 40454 55681
rect 40396 55641 40408 55675
rect 40442 55672 40454 55675
rect 40494 55672 40500 55684
rect 40442 55644 40500 55672
rect 40442 55641 40454 55644
rect 40396 55635 40454 55641
rect 40494 55632 40500 55644
rect 40552 55632 40558 55684
rect 46584 55672 46612 55768
rect 46845 55743 46903 55749
rect 46845 55709 46857 55743
rect 46891 55740 46903 55743
rect 46934 55740 46940 55752
rect 46891 55712 46940 55740
rect 46891 55709 46903 55712
rect 46845 55703 46903 55709
rect 46934 55700 46940 55712
rect 46992 55700 46998 55752
rect 47581 55743 47639 55749
rect 47581 55709 47593 55743
rect 47627 55740 47639 55743
rect 48516 55740 48544 55780
rect 50157 55777 50169 55780
rect 50203 55808 50215 55811
rect 50522 55808 50528 55820
rect 50203 55780 50528 55808
rect 50203 55777 50215 55780
rect 50157 55771 50215 55777
rect 50522 55768 50528 55780
rect 50580 55768 50586 55820
rect 47627 55712 48544 55740
rect 47627 55709 47639 55712
rect 47581 55703 47639 55709
rect 48590 55700 48596 55752
rect 48648 55740 48654 55752
rect 50338 55740 50344 55752
rect 48648 55712 48693 55740
rect 50299 55712 50344 55740
rect 48648 55700 48654 55712
rect 50338 55700 50344 55712
rect 50396 55700 50402 55752
rect 47857 55675 47915 55681
rect 47857 55672 47869 55675
rect 46584 55644 47869 55672
rect 47857 55641 47869 55644
rect 47903 55641 47915 55675
rect 47857 55635 47915 55641
rect 41509 55607 41567 55613
rect 41509 55604 41521 55607
rect 39592 55576 41521 55604
rect 41509 55573 41521 55576
rect 41555 55573 41567 55607
rect 41509 55567 41567 55573
rect 47581 55607 47639 55613
rect 47581 55573 47593 55607
rect 47627 55604 47639 55607
rect 47946 55604 47952 55616
rect 47627 55576 47952 55604
rect 47627 55573 47639 55576
rect 47581 55567 47639 55573
rect 47946 55564 47952 55576
rect 48004 55564 48010 55616
rect 1104 55514 68816 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 68816 55514
rect 1104 55440 68816 55462
rect 25406 55400 25412 55412
rect 25367 55372 25412 55400
rect 25406 55360 25412 55372
rect 25464 55360 25470 55412
rect 27154 55360 27160 55412
rect 27212 55400 27218 55412
rect 27709 55403 27767 55409
rect 27709 55400 27721 55403
rect 27212 55372 27721 55400
rect 27212 55360 27218 55372
rect 27709 55369 27721 55372
rect 27755 55369 27767 55403
rect 28534 55400 28540 55412
rect 28495 55372 28540 55400
rect 27709 55363 27767 55369
rect 28534 55360 28540 55372
rect 28592 55360 28598 55412
rect 31386 55400 31392 55412
rect 31347 55372 31392 55400
rect 31386 55360 31392 55372
rect 31444 55360 31450 55412
rect 32674 55400 32680 55412
rect 32635 55372 32680 55400
rect 32674 55360 32680 55372
rect 32732 55360 32738 55412
rect 36630 55400 36636 55412
rect 36591 55372 36636 55400
rect 36630 55360 36636 55372
rect 36688 55360 36694 55412
rect 39022 55360 39028 55412
rect 39080 55360 39086 55412
rect 40494 55400 40500 55412
rect 40455 55372 40500 55400
rect 40494 55360 40500 55372
rect 40552 55360 40558 55412
rect 43898 55400 43904 55412
rect 43859 55372 43904 55400
rect 43898 55360 43904 55372
rect 43956 55360 43962 55412
rect 47578 55400 47584 55412
rect 47539 55372 47584 55400
rect 47578 55360 47584 55372
rect 47636 55360 47642 55412
rect 14452 55335 14510 55341
rect 14452 55301 14464 55335
rect 14498 55332 14510 55335
rect 14642 55332 14648 55344
rect 14498 55304 14648 55332
rect 14498 55301 14510 55304
rect 14452 55295 14510 55301
rect 14642 55292 14648 55304
rect 14700 55292 14706 55344
rect 36262 55332 36268 55344
rect 35820 55304 36268 55332
rect 13633 55267 13691 55273
rect 13633 55233 13645 55267
rect 13679 55264 13691 55267
rect 13814 55264 13820 55276
rect 13679 55236 13820 55264
rect 13679 55233 13691 55236
rect 13633 55227 13691 55233
rect 13814 55224 13820 55236
rect 13872 55224 13878 55276
rect 16942 55264 16948 55276
rect 16903 55236 16948 55264
rect 16942 55224 16948 55236
rect 17000 55224 17006 55276
rect 17212 55267 17270 55273
rect 17212 55233 17224 55267
rect 17258 55264 17270 55267
rect 17678 55264 17684 55276
rect 17258 55236 17684 55264
rect 17258 55233 17270 55236
rect 17212 55227 17270 55233
rect 17678 55224 17684 55236
rect 17736 55224 17742 55276
rect 18230 55224 18236 55276
rect 18288 55264 18294 55276
rect 18969 55267 19027 55273
rect 18969 55264 18981 55267
rect 18288 55236 18981 55264
rect 18288 55224 18294 55236
rect 18969 55233 18981 55236
rect 19015 55233 19027 55267
rect 18969 55227 19027 55233
rect 22922 55224 22928 55276
rect 22980 55264 22986 55276
rect 23293 55267 23351 55273
rect 23293 55264 23305 55267
rect 22980 55236 23305 55264
rect 22980 55224 22986 55236
rect 23293 55233 23305 55236
rect 23339 55233 23351 55267
rect 25130 55264 25136 55276
rect 25091 55236 25136 55264
rect 23293 55227 23351 55233
rect 25130 55224 25136 55236
rect 25188 55224 25194 55276
rect 25225 55267 25283 55273
rect 25225 55233 25237 55267
rect 25271 55264 25283 55267
rect 25498 55264 25504 55276
rect 25271 55236 25504 55264
rect 25271 55233 25283 55236
rect 25225 55227 25283 55233
rect 25498 55224 25504 55236
rect 25556 55224 25562 55276
rect 25682 55264 25688 55276
rect 25608 55236 25688 55264
rect 13725 55199 13783 55205
rect 13725 55165 13737 55199
rect 13771 55196 13783 55199
rect 14185 55199 14243 55205
rect 14185 55196 14197 55199
rect 13771 55168 14197 55196
rect 13771 55165 13783 55168
rect 13725 55159 13783 55165
rect 14185 55165 14197 55168
rect 14231 55165 14243 55199
rect 18785 55199 18843 55205
rect 18785 55196 18797 55199
rect 14185 55159 14243 55165
rect 18340 55168 18797 55196
rect 15562 55060 15568 55072
rect 15523 55032 15568 55060
rect 15562 55020 15568 55032
rect 15620 55020 15626 55072
rect 18046 55020 18052 55072
rect 18104 55060 18110 55072
rect 18340 55069 18368 55168
rect 18785 55165 18797 55168
rect 18831 55165 18843 55199
rect 18785 55159 18843 55165
rect 23569 55199 23627 55205
rect 23569 55165 23581 55199
rect 23615 55196 23627 55199
rect 25608 55196 25636 55236
rect 25682 55224 25688 55236
rect 25740 55264 25746 55276
rect 27617 55267 27675 55273
rect 27617 55264 27629 55267
rect 25740 55236 27629 55264
rect 25740 55224 25746 55236
rect 27617 55233 27629 55236
rect 27663 55233 27675 55267
rect 28718 55264 28724 55276
rect 28679 55236 28724 55264
rect 27617 55227 27675 55233
rect 28718 55224 28724 55236
rect 28776 55224 28782 55276
rect 30742 55224 30748 55276
rect 30800 55264 30806 55276
rect 31573 55267 31631 55273
rect 31573 55264 31585 55267
rect 30800 55236 31585 55264
rect 30800 55224 30806 55236
rect 31573 55233 31585 55236
rect 31619 55233 31631 55267
rect 31573 55227 31631 55233
rect 32214 55224 32220 55276
rect 32272 55264 32278 55276
rect 32490 55264 32496 55276
rect 32272 55236 32496 55264
rect 32272 55224 32278 55236
rect 32490 55224 32496 55236
rect 32548 55264 32554 55276
rect 32585 55267 32643 55273
rect 32585 55264 32597 55267
rect 32548 55236 32597 55264
rect 32548 55224 32554 55236
rect 32585 55233 32597 55236
rect 32631 55233 32643 55267
rect 32585 55227 32643 55233
rect 33042 55224 33048 55276
rect 33100 55264 33106 55276
rect 33597 55267 33655 55273
rect 33597 55264 33609 55267
rect 33100 55236 33609 55264
rect 33100 55224 33106 55236
rect 33597 55233 33609 55236
rect 33643 55233 33655 55267
rect 33597 55227 33655 55233
rect 33864 55267 33922 55273
rect 33864 55233 33876 55267
rect 33910 55264 33922 55267
rect 34698 55264 34704 55276
rect 33910 55236 34704 55264
rect 33910 55233 33922 55236
rect 33864 55227 33922 55233
rect 34698 55224 34704 55236
rect 34756 55224 34762 55276
rect 35526 55224 35532 55276
rect 35584 55264 35590 55276
rect 35820 55273 35848 55304
rect 36262 55292 36268 55304
rect 36320 55292 36326 55344
rect 36722 55292 36728 55344
rect 36780 55332 36786 55344
rect 37737 55335 37795 55341
rect 37737 55332 37749 55335
rect 36780 55304 37749 55332
rect 36780 55292 36786 55304
rect 37737 55301 37749 55304
rect 37783 55301 37795 55335
rect 39040 55332 39068 55360
rect 37737 55295 37795 55301
rect 38948 55304 39068 55332
rect 45848 55304 50384 55332
rect 35805 55267 35863 55273
rect 35805 55264 35817 55267
rect 35584 55236 35817 55264
rect 35584 55224 35590 55236
rect 35805 55233 35817 55236
rect 35851 55233 35863 55267
rect 35805 55227 35863 55233
rect 35989 55267 36047 55273
rect 35989 55233 36001 55267
rect 36035 55264 36047 55267
rect 36078 55264 36084 55276
rect 36035 55236 36084 55264
rect 36035 55233 36047 55236
rect 35989 55227 36047 55233
rect 36078 55224 36084 55236
rect 36136 55224 36142 55276
rect 36541 55267 36599 55273
rect 36541 55233 36553 55267
rect 36587 55264 36599 55267
rect 37182 55264 37188 55276
rect 36587 55236 37188 55264
rect 36587 55233 36599 55236
rect 36541 55227 36599 55233
rect 37182 55224 37188 55236
rect 37240 55224 37246 55276
rect 38948 55273 38976 55304
rect 45848 55276 45876 55304
rect 38933 55267 38991 55273
rect 38933 55233 38945 55267
rect 38979 55233 38991 55267
rect 39114 55264 39120 55276
rect 39075 55236 39120 55264
rect 38933 55227 38991 55233
rect 39114 55224 39120 55236
rect 39172 55224 39178 55276
rect 40681 55267 40739 55273
rect 40681 55233 40693 55267
rect 40727 55264 40739 55267
rect 41322 55264 41328 55276
rect 40727 55236 41328 55264
rect 40727 55233 40739 55236
rect 40681 55227 40739 55233
rect 41322 55224 41328 55236
rect 41380 55224 41386 55276
rect 42518 55264 42524 55276
rect 42479 55236 42524 55264
rect 42518 55224 42524 55236
rect 42576 55224 42582 55276
rect 42788 55267 42846 55273
rect 42788 55233 42800 55267
rect 42834 55264 42846 55267
rect 43162 55264 43168 55276
rect 42834 55236 43168 55264
rect 42834 55233 42846 55236
rect 42788 55227 42846 55233
rect 43162 55224 43168 55236
rect 43220 55224 43226 55276
rect 45830 55264 45836 55276
rect 45791 55236 45836 55264
rect 45830 55224 45836 55236
rect 45888 55224 45894 55276
rect 47762 55264 47768 55276
rect 47723 55236 47768 55264
rect 47762 55224 47768 55236
rect 47820 55224 47826 55276
rect 48498 55264 48504 55276
rect 48459 55236 48504 55264
rect 48498 55224 48504 55236
rect 48556 55224 48562 55276
rect 50356 55273 50384 55304
rect 50341 55267 50399 55273
rect 50341 55233 50353 55267
rect 50387 55233 50399 55267
rect 51258 55264 51264 55276
rect 51219 55236 51264 55264
rect 50341 55227 50399 55233
rect 51258 55224 51264 55236
rect 51316 55224 51322 55276
rect 23615 55168 25636 55196
rect 23615 55165 23627 55168
rect 23569 55159 23627 55165
rect 39022 55156 39028 55208
rect 39080 55196 39086 55208
rect 39209 55199 39267 55205
rect 39209 55196 39221 55199
rect 39080 55168 39221 55196
rect 39080 55156 39086 55168
rect 39209 55165 39221 55168
rect 39255 55165 39267 55199
rect 39209 55159 39267 55165
rect 40957 55199 41015 55205
rect 40957 55165 40969 55199
rect 41003 55196 41015 55199
rect 42426 55196 42432 55208
rect 41003 55168 42432 55196
rect 41003 55165 41015 55168
rect 40957 55159 41015 55165
rect 42426 55156 42432 55168
rect 42484 55156 42490 55208
rect 35986 55088 35992 55140
rect 36044 55128 36050 55140
rect 36262 55128 36268 55140
rect 36044 55100 36268 55128
rect 36044 55088 36050 55100
rect 36262 55088 36268 55100
rect 36320 55088 36326 55140
rect 38749 55131 38807 55137
rect 38749 55097 38761 55131
rect 38795 55128 38807 55131
rect 40865 55131 40923 55137
rect 40865 55128 40877 55131
rect 38795 55100 40877 55128
rect 38795 55097 38807 55100
rect 38749 55091 38807 55097
rect 40865 55097 40877 55100
rect 40911 55097 40923 55131
rect 40865 55091 40923 55097
rect 18325 55063 18383 55069
rect 18325 55060 18337 55063
rect 18104 55032 18337 55060
rect 18104 55020 18110 55032
rect 18325 55029 18337 55032
rect 18371 55029 18383 55063
rect 19150 55060 19156 55072
rect 19111 55032 19156 55060
rect 18325 55023 18383 55029
rect 19150 55020 19156 55032
rect 19208 55020 19214 55072
rect 34977 55063 35035 55069
rect 34977 55029 34989 55063
rect 35023 55060 35035 55063
rect 35434 55060 35440 55072
rect 35023 55032 35440 55060
rect 35023 55029 35035 55032
rect 34977 55023 35035 55029
rect 35434 55020 35440 55032
rect 35492 55020 35498 55072
rect 35802 55060 35808 55072
rect 35763 55032 35808 55060
rect 35802 55020 35808 55032
rect 35860 55020 35866 55072
rect 37826 55060 37832 55072
rect 37787 55032 37832 55060
rect 37826 55020 37832 55032
rect 37884 55020 37890 55072
rect 45738 55060 45744 55072
rect 45699 55032 45744 55060
rect 45738 55020 45744 55032
rect 45796 55020 45802 55072
rect 48314 55060 48320 55072
rect 48275 55032 48320 55060
rect 48314 55020 48320 55032
rect 48372 55020 48378 55072
rect 50341 55063 50399 55069
rect 50341 55029 50353 55063
rect 50387 55060 50399 55063
rect 50430 55060 50436 55072
rect 50387 55032 50436 55060
rect 50387 55029 50399 55032
rect 50341 55023 50399 55029
rect 50430 55020 50436 55032
rect 50488 55020 50494 55072
rect 51074 55060 51080 55072
rect 51035 55032 51080 55060
rect 51074 55020 51080 55032
rect 51132 55020 51138 55072
rect 1104 54970 68816 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 65654 54970
rect 65706 54918 65718 54970
rect 65770 54918 65782 54970
rect 65834 54918 65846 54970
rect 65898 54918 65910 54970
rect 65962 54918 68816 54970
rect 1104 54896 68816 54918
rect 15286 54856 15292 54868
rect 15247 54828 15292 54856
rect 15286 54816 15292 54828
rect 15344 54816 15350 54868
rect 17678 54856 17684 54868
rect 17639 54828 17684 54856
rect 17678 54816 17684 54828
rect 17736 54816 17742 54868
rect 21729 54859 21787 54865
rect 21729 54825 21741 54859
rect 21775 54856 21787 54859
rect 22186 54856 22192 54868
rect 21775 54828 22192 54856
rect 21775 54825 21787 54828
rect 21729 54819 21787 54825
rect 22186 54816 22192 54828
rect 22244 54816 22250 54868
rect 34698 54856 34704 54868
rect 34659 54828 34704 54856
rect 34698 54816 34704 54828
rect 34756 54816 34762 54868
rect 35069 54859 35127 54865
rect 35069 54825 35081 54859
rect 35115 54856 35127 54859
rect 35710 54856 35716 54868
rect 35115 54828 35716 54856
rect 35115 54825 35127 54828
rect 35069 54819 35127 54825
rect 35710 54816 35716 54828
rect 35768 54856 35774 54868
rect 38654 54856 38660 54868
rect 35768 54828 35940 54856
rect 38615 54828 38660 54856
rect 35768 54816 35774 54828
rect 20809 54791 20867 54797
rect 20809 54757 20821 54791
rect 20855 54788 20867 54791
rect 21818 54788 21824 54800
rect 20855 54760 21824 54788
rect 20855 54757 20867 54760
rect 20809 54751 20867 54757
rect 21818 54748 21824 54760
rect 21876 54748 21882 54800
rect 22830 54788 22836 54800
rect 22020 54760 22836 54788
rect 21726 54720 21732 54732
rect 21008 54692 21732 54720
rect 15013 54655 15071 54661
rect 15013 54621 15025 54655
rect 15059 54621 15071 54655
rect 15013 54615 15071 54621
rect 15105 54655 15163 54661
rect 15105 54621 15117 54655
rect 15151 54652 15163 54655
rect 15194 54652 15200 54664
rect 15151 54624 15200 54652
rect 15151 54621 15163 54624
rect 15105 54615 15163 54621
rect 15028 54584 15056 54615
rect 15194 54612 15200 54624
rect 15252 54612 15258 54664
rect 17865 54655 17923 54661
rect 17865 54621 17877 54655
rect 17911 54652 17923 54655
rect 19150 54652 19156 54664
rect 17911 54624 19156 54652
rect 17911 54621 17923 54624
rect 17865 54615 17923 54621
rect 19150 54612 19156 54624
rect 19208 54612 19214 54664
rect 19613 54655 19671 54661
rect 19613 54621 19625 54655
rect 19659 54652 19671 54655
rect 19978 54652 19984 54664
rect 19659 54624 19984 54652
rect 19659 54621 19671 54624
rect 19613 54615 19671 54621
rect 19978 54612 19984 54624
rect 20036 54612 20042 54664
rect 20346 54652 20352 54664
rect 20307 54624 20352 54652
rect 20346 54612 20352 54624
rect 20404 54612 20410 54664
rect 21008 54661 21036 54692
rect 21726 54680 21732 54692
rect 21784 54680 21790 54732
rect 22020 54661 22048 54760
rect 22830 54748 22836 54760
rect 22888 54748 22894 54800
rect 31389 54791 31447 54797
rect 31389 54757 31401 54791
rect 31435 54788 31447 54791
rect 33318 54788 33324 54800
rect 31435 54760 33324 54788
rect 31435 54757 31447 54760
rect 31389 54751 31447 54757
rect 33318 54748 33324 54760
rect 33376 54748 33382 54800
rect 35621 54791 35679 54797
rect 35621 54757 35633 54791
rect 35667 54757 35679 54791
rect 35621 54751 35679 54757
rect 24026 54720 24032 54732
rect 22112 54692 24032 54720
rect 22112 54661 22140 54692
rect 20993 54655 21051 54661
rect 20993 54621 21005 54655
rect 21039 54621 21051 54655
rect 21269 54655 21327 54661
rect 21269 54652 21281 54655
rect 20993 54615 21051 54621
rect 21100 54624 21281 54652
rect 15562 54584 15568 54596
rect 15028 54556 15568 54584
rect 15562 54544 15568 54556
rect 15620 54584 15626 54596
rect 18230 54584 18236 54596
rect 15620 54556 18236 54584
rect 15620 54544 15626 54556
rect 18230 54544 18236 54556
rect 18288 54544 18294 54596
rect 19242 54544 19248 54596
rect 19300 54584 19306 54596
rect 21100 54584 21128 54624
rect 21269 54621 21281 54624
rect 21315 54621 21327 54655
rect 21269 54615 21327 54621
rect 22005 54655 22063 54661
rect 22005 54621 22017 54655
rect 22051 54621 22063 54655
rect 22005 54615 22063 54621
rect 22097 54655 22155 54661
rect 22097 54621 22109 54655
rect 22143 54621 22155 54655
rect 22097 54615 22155 54621
rect 22189 54655 22247 54661
rect 22189 54621 22201 54655
rect 22235 54621 22247 54655
rect 22189 54615 22247 54621
rect 22373 54655 22431 54661
rect 22373 54621 22385 54655
rect 22419 54621 22431 54655
rect 22373 54615 22431 54621
rect 19300 54556 21128 54584
rect 21177 54587 21235 54593
rect 19300 54544 19306 54556
rect 21177 54553 21189 54587
rect 21223 54584 21235 54587
rect 21223 54556 21864 54584
rect 21223 54553 21235 54556
rect 21177 54547 21235 54553
rect 17494 54476 17500 54528
rect 17552 54516 17558 54528
rect 19334 54516 19340 54528
rect 17552 54488 19340 54516
rect 17552 54476 17558 54488
rect 19334 54476 19340 54488
rect 19392 54476 19398 54528
rect 19426 54476 19432 54528
rect 19484 54516 19490 54528
rect 19613 54519 19671 54525
rect 19613 54516 19625 54519
rect 19484 54488 19625 54516
rect 19484 54476 19490 54488
rect 19613 54485 19625 54488
rect 19659 54485 19671 54519
rect 20162 54516 20168 54528
rect 20123 54488 20168 54516
rect 19613 54479 19671 54485
rect 20162 54476 20168 54488
rect 20220 54476 20226 54528
rect 21836 54516 21864 54556
rect 21910 54544 21916 54596
rect 21968 54584 21974 54596
rect 22204 54584 22232 54615
rect 21968 54556 22232 54584
rect 22388 54584 22416 54615
rect 22830 54612 22836 54664
rect 22888 54652 22894 54664
rect 23308 54661 23336 54692
rect 24026 54680 24032 54692
rect 24084 54680 24090 54732
rect 31662 54720 31668 54732
rect 31575 54692 31668 54720
rect 23201 54655 23259 54661
rect 23201 54652 23213 54655
rect 22888 54624 23213 54652
rect 22888 54612 22894 54624
rect 23201 54621 23213 54624
rect 23247 54621 23259 54655
rect 23201 54615 23259 54621
rect 23293 54655 23351 54661
rect 23293 54621 23305 54655
rect 23339 54621 23351 54655
rect 23293 54615 23351 54621
rect 23382 54612 23388 54664
rect 23440 54652 23446 54664
rect 23569 54655 23627 54661
rect 23440 54624 23485 54652
rect 23440 54612 23446 54624
rect 23569 54621 23581 54655
rect 23615 54621 23627 54655
rect 25406 54652 25412 54664
rect 25367 54624 25412 54652
rect 23569 54615 23627 54621
rect 23014 54584 23020 54596
rect 22388 54556 23020 54584
rect 21968 54544 21974 54556
rect 23014 54544 23020 54556
rect 23072 54584 23078 54596
rect 23584 54584 23612 54615
rect 25406 54612 25412 54624
rect 25464 54612 25470 54664
rect 28994 54652 29000 54664
rect 28955 54624 29000 54652
rect 28994 54612 29000 54624
rect 29052 54612 29058 54664
rect 30101 54655 30159 54661
rect 30101 54621 30113 54655
rect 30147 54652 30159 54655
rect 30558 54652 30564 54664
rect 30147 54624 30564 54652
rect 30147 54621 30159 54624
rect 30101 54615 30159 54621
rect 30558 54612 30564 54624
rect 30616 54612 30622 54664
rect 31588 54661 31616 54692
rect 31662 54680 31668 54692
rect 31720 54720 31726 54732
rect 32585 54723 32643 54729
rect 32585 54720 32597 54723
rect 31720 54692 32597 54720
rect 31720 54680 31726 54692
rect 32585 54689 32597 54692
rect 32631 54689 32643 54723
rect 35636 54720 35664 54751
rect 32585 54683 32643 54689
rect 34900 54692 35664 54720
rect 31573 54655 31631 54661
rect 31573 54621 31585 54655
rect 31619 54621 31631 54655
rect 31754 54652 31760 54664
rect 31715 54624 31760 54652
rect 31573 54615 31631 54621
rect 31754 54612 31760 54624
rect 31812 54612 31818 54664
rect 31846 54612 31852 54664
rect 31904 54652 31910 54664
rect 34900 54661 34928 54692
rect 34885 54655 34943 54661
rect 31904 54624 31949 54652
rect 31904 54612 31910 54624
rect 34885 54621 34897 54655
rect 34931 54621 34943 54655
rect 34885 54615 34943 54621
rect 35161 54655 35219 54661
rect 35161 54621 35173 54655
rect 35207 54652 35219 54655
rect 35434 54652 35440 54664
rect 35207 54624 35440 54652
rect 35207 54621 35219 54624
rect 35161 54615 35219 54621
rect 35434 54612 35440 54624
rect 35492 54652 35498 54664
rect 35710 54652 35716 54664
rect 35492 54624 35716 54652
rect 35492 54612 35498 54624
rect 35710 54612 35716 54624
rect 35768 54652 35774 54664
rect 35912 54661 35940 54828
rect 38654 54816 38660 54828
rect 38712 54816 38718 54868
rect 45189 54859 45247 54865
rect 45189 54825 45201 54859
rect 45235 54856 45247 54859
rect 45370 54856 45376 54868
rect 45235 54828 45376 54856
rect 45235 54825 45247 54828
rect 45189 54819 45247 54825
rect 41322 54720 41328 54732
rect 38488 54692 41328 54720
rect 38488 54661 38516 54692
rect 41322 54680 41328 54692
rect 41380 54680 41386 54732
rect 45204 54720 45232 54819
rect 45370 54816 45376 54828
rect 45428 54856 45434 54868
rect 46934 54856 46940 54868
rect 45428 54828 46940 54856
rect 45428 54816 45434 54828
rect 46934 54816 46940 54828
rect 46992 54816 46998 54868
rect 45738 54720 45744 54732
rect 44192 54692 45232 54720
rect 45699 54692 45744 54720
rect 35805 54655 35863 54661
rect 35805 54652 35817 54655
rect 35768 54624 35817 54652
rect 35768 54612 35774 54624
rect 35805 54621 35817 54624
rect 35851 54621 35863 54655
rect 35805 54615 35863 54621
rect 35897 54655 35955 54661
rect 35897 54621 35909 54655
rect 35943 54621 35955 54655
rect 35897 54615 35955 54621
rect 38473 54655 38531 54661
rect 38473 54621 38485 54655
rect 38519 54621 38531 54655
rect 38473 54615 38531 54621
rect 38749 54655 38807 54661
rect 38749 54621 38761 54655
rect 38795 54652 38807 54655
rect 38930 54652 38936 54664
rect 38795 54624 38936 54652
rect 38795 54621 38807 54624
rect 38749 54615 38807 54621
rect 38930 54612 38936 54624
rect 38988 54612 38994 54664
rect 42981 54655 43039 54661
rect 42981 54621 42993 54655
rect 43027 54652 43039 54655
rect 43070 54652 43076 54664
rect 43027 54624 43076 54652
rect 43027 54621 43039 54624
rect 42981 54615 43039 54621
rect 43070 54612 43076 54624
rect 43128 54612 43134 54664
rect 44192 54661 44220 54692
rect 45738 54680 45744 54692
rect 45796 54680 45802 54732
rect 50430 54720 50436 54732
rect 50391 54692 50436 54720
rect 50430 54680 50436 54692
rect 50488 54680 50494 54732
rect 44177 54655 44235 54661
rect 44177 54621 44189 54655
rect 44223 54621 44235 54655
rect 45002 54652 45008 54664
rect 44963 54624 45008 54652
rect 44177 54615 44235 54621
rect 45002 54612 45008 54624
rect 45060 54612 45066 54664
rect 47670 54652 47676 54664
rect 47631 54624 47676 54652
rect 47670 54612 47676 54624
rect 47728 54612 47734 54664
rect 47940 54655 47998 54661
rect 47940 54621 47952 54655
rect 47986 54652 47998 54655
rect 48314 54652 48320 54664
rect 47986 54624 48320 54652
rect 47986 54621 47998 54624
rect 47940 54615 47998 54621
rect 48314 54612 48320 54624
rect 48372 54612 48378 54664
rect 50700 54655 50758 54661
rect 50700 54621 50712 54655
rect 50746 54652 50758 54655
rect 51074 54652 51080 54664
rect 50746 54624 51080 54652
rect 50746 54621 50758 54624
rect 50700 54615 50758 54621
rect 51074 54612 51080 54624
rect 51132 54612 51138 54664
rect 23072 54556 23612 54584
rect 28813 54587 28871 54593
rect 23072 54544 23078 54556
rect 28813 54553 28825 54587
rect 28859 54584 28871 54587
rect 30006 54584 30012 54596
rect 28859 54556 30012 54584
rect 28859 54553 28871 54556
rect 28813 54547 28871 54553
rect 30006 54544 30012 54556
rect 30064 54544 30070 54596
rect 32398 54584 32404 54596
rect 32311 54556 32404 54584
rect 32398 54544 32404 54556
rect 32456 54584 32462 54596
rect 35621 54587 35679 54593
rect 32456 54556 33180 54584
rect 32456 54544 32462 54556
rect 22278 54516 22284 54528
rect 21836 54488 22284 54516
rect 22278 54476 22284 54488
rect 22336 54476 22342 54528
rect 22925 54519 22983 54525
rect 22925 54485 22937 54519
rect 22971 54516 22983 54519
rect 23290 54516 23296 54528
rect 22971 54488 23296 54516
rect 22971 54485 22983 54488
rect 22925 54479 22983 54485
rect 23290 54476 23296 54488
rect 23348 54476 23354 54528
rect 25130 54476 25136 54528
rect 25188 54516 25194 54528
rect 25225 54519 25283 54525
rect 25225 54516 25237 54519
rect 25188 54488 25237 54516
rect 25188 54476 25194 54488
rect 25225 54485 25237 54488
rect 25271 54485 25283 54519
rect 25225 54479 25283 54485
rect 29822 54476 29828 54528
rect 29880 54516 29886 54528
rect 30101 54519 30159 54525
rect 30101 54516 30113 54519
rect 29880 54488 30113 54516
rect 29880 54476 29886 54488
rect 30101 54485 30113 54488
rect 30147 54485 30159 54519
rect 33152 54516 33180 54556
rect 35621 54553 35633 54587
rect 35667 54584 35679 54587
rect 36722 54584 36728 54596
rect 35667 54556 36728 54584
rect 35667 54553 35679 54556
rect 35621 54547 35679 54553
rect 36722 54544 36728 54556
rect 36780 54584 36786 54596
rect 41414 54584 41420 54596
rect 36780 54556 41420 54584
rect 36780 54544 36786 54556
rect 41414 54544 41420 54556
rect 41472 54584 41478 54596
rect 41598 54584 41604 54596
rect 41472 54556 41604 54584
rect 41472 54544 41478 54556
rect 41598 54544 41604 54556
rect 41656 54544 41662 54596
rect 43162 54584 43168 54596
rect 43123 54556 43168 54584
rect 43162 54544 43168 54556
rect 43220 54544 43226 54596
rect 45646 54544 45652 54596
rect 45704 54584 45710 54596
rect 45986 54587 46044 54593
rect 45986 54584 45998 54587
rect 45704 54556 45998 54584
rect 45704 54544 45710 54556
rect 45986 54553 45998 54556
rect 46032 54553 46044 54587
rect 45986 54547 46044 54553
rect 38102 54516 38108 54528
rect 33152 54488 38108 54516
rect 30101 54479 30159 54485
rect 38102 54476 38108 54488
rect 38160 54476 38166 54528
rect 38286 54516 38292 54528
rect 38247 54488 38292 54516
rect 38286 54476 38292 54488
rect 38344 54476 38350 54528
rect 43622 54476 43628 54528
rect 43680 54516 43686 54528
rect 44269 54519 44327 54525
rect 44269 54516 44281 54519
rect 43680 54488 44281 54516
rect 43680 54476 43686 54488
rect 44269 54485 44281 54488
rect 44315 54485 44327 54519
rect 44269 54479 44327 54485
rect 46566 54476 46572 54528
rect 46624 54516 46630 54528
rect 47121 54519 47179 54525
rect 47121 54516 47133 54519
rect 46624 54488 47133 54516
rect 46624 54476 46630 54488
rect 47121 54485 47133 54488
rect 47167 54485 47179 54519
rect 47121 54479 47179 54485
rect 48682 54476 48688 54528
rect 48740 54516 48746 54528
rect 49053 54519 49111 54525
rect 49053 54516 49065 54519
rect 48740 54488 49065 54516
rect 48740 54476 48746 54488
rect 49053 54485 49065 54488
rect 49099 54485 49111 54519
rect 49053 54479 49111 54485
rect 49878 54476 49884 54528
rect 49936 54516 49942 54528
rect 51813 54519 51871 54525
rect 51813 54516 51825 54519
rect 49936 54488 51825 54516
rect 49936 54476 49942 54488
rect 51813 54485 51825 54488
rect 51859 54485 51871 54519
rect 51813 54479 51871 54485
rect 1104 54426 68816 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 68816 54426
rect 1104 54352 68816 54374
rect 33134 54312 33140 54324
rect 6380 54284 33140 54312
rect 6380 54185 6408 54284
rect 33134 54272 33140 54284
rect 33192 54312 33198 54324
rect 33505 54315 33563 54321
rect 33505 54312 33517 54315
rect 33192 54284 33517 54312
rect 33192 54272 33198 54284
rect 33505 54281 33517 54284
rect 33551 54281 33563 54315
rect 45186 54312 45192 54324
rect 33505 54275 33563 54281
rect 41386 54284 45192 54312
rect 19153 54247 19211 54253
rect 19153 54213 19165 54247
rect 19199 54244 19211 54247
rect 19242 54244 19248 54256
rect 19199 54216 19248 54244
rect 19199 54213 19211 54216
rect 19153 54207 19211 54213
rect 19242 54204 19248 54216
rect 19300 54204 19306 54256
rect 19880 54247 19938 54253
rect 19880 54213 19892 54247
rect 19926 54244 19938 54247
rect 20162 54244 20168 54256
rect 19926 54216 20168 54244
rect 19926 54213 19938 54216
rect 19880 54207 19938 54213
rect 20162 54204 20168 54216
rect 20220 54204 20226 54256
rect 21821 54247 21879 54253
rect 21821 54213 21833 54247
rect 21867 54244 21879 54247
rect 21910 54244 21916 54256
rect 21867 54216 21916 54244
rect 21867 54213 21879 54216
rect 21821 54207 21879 54213
rect 21910 54204 21916 54216
rect 21968 54204 21974 54256
rect 22186 54244 22192 54256
rect 22147 54216 22192 54244
rect 22186 54204 22192 54216
rect 22244 54204 22250 54256
rect 28994 54244 29000 54256
rect 23124 54216 29000 54244
rect 6365 54179 6423 54185
rect 6365 54145 6377 54179
rect 6411 54145 6423 54179
rect 6365 54139 6423 54145
rect 15933 54179 15991 54185
rect 15933 54145 15945 54179
rect 15979 54176 15991 54179
rect 16574 54176 16580 54188
rect 15979 54148 16580 54176
rect 15979 54145 15991 54148
rect 15933 54139 15991 54145
rect 16574 54136 16580 54148
rect 16632 54136 16638 54188
rect 17313 54179 17371 54185
rect 17313 54145 17325 54179
rect 17359 54176 17371 54179
rect 17359 54148 17724 54176
rect 17359 54145 17371 54148
rect 17313 54139 17371 54145
rect 6546 54108 6552 54120
rect 6507 54080 6552 54108
rect 6546 54068 6552 54080
rect 6604 54068 6610 54120
rect 6917 54111 6975 54117
rect 6917 54077 6929 54111
rect 6963 54077 6975 54111
rect 6917 54071 6975 54077
rect 15749 54111 15807 54117
rect 15749 54077 15761 54111
rect 15795 54108 15807 54111
rect 17494 54108 17500 54120
rect 15795 54080 16988 54108
rect 17455 54080 17500 54108
rect 15795 54077 15807 54080
rect 15749 54071 15807 54077
rect 3510 54000 3516 54052
rect 3568 54040 3574 54052
rect 6932 54040 6960 54071
rect 3568 54012 6960 54040
rect 3568 54000 3574 54012
rect 16960 53984 16988 54080
rect 17494 54068 17500 54080
rect 17552 54068 17558 54120
rect 17696 54108 17724 54148
rect 18230 54136 18236 54188
rect 18288 54176 18294 54188
rect 18288 54148 18333 54176
rect 18288 54136 18294 54148
rect 19426 54136 19432 54188
rect 19484 54176 19490 54188
rect 19613 54179 19671 54185
rect 19613 54176 19625 54179
rect 19484 54148 19625 54176
rect 19484 54136 19490 54148
rect 19613 54145 19625 54148
rect 19659 54145 19671 54179
rect 19613 54139 19671 54145
rect 21726 54136 21732 54188
rect 21784 54176 21790 54188
rect 22005 54179 22063 54185
rect 22005 54176 22017 54179
rect 21784 54148 22017 54176
rect 21784 54136 21790 54148
rect 22005 54145 22017 54148
rect 22051 54145 22063 54179
rect 22005 54139 22063 54145
rect 22281 54179 22339 54185
rect 22281 54145 22293 54179
rect 22327 54145 22339 54179
rect 23124 54176 23152 54216
rect 28994 54204 29000 54216
rect 29052 54244 29058 54256
rect 37820 54247 37878 54253
rect 29052 54216 31754 54244
rect 29052 54204 29058 54216
rect 23198 54176 23204 54188
rect 23124 54148 23204 54176
rect 22281 54139 22339 54145
rect 18046 54108 18052 54120
rect 17696 54080 18052 54108
rect 18046 54068 18052 54080
rect 18104 54068 18110 54120
rect 18322 54068 18328 54120
rect 18380 54117 18386 54120
rect 18380 54111 18408 54117
rect 18396 54077 18408 54111
rect 18380 54071 18408 54077
rect 18380 54068 18386 54071
rect 18506 54068 18512 54120
rect 18564 54108 18570 54120
rect 18564 54080 18609 54108
rect 18564 54068 18570 54080
rect 20622 54068 20628 54120
rect 20680 54108 20686 54120
rect 22296 54108 22324 54139
rect 23198 54136 23204 54148
rect 23256 54136 23262 54188
rect 23290 54136 23296 54188
rect 23348 54176 23354 54188
rect 23457 54179 23515 54185
rect 23457 54176 23469 54179
rect 23348 54148 23469 54176
rect 23348 54136 23354 54148
rect 23457 54145 23469 54148
rect 23503 54145 23515 54179
rect 23457 54139 23515 54145
rect 24946 54136 24952 54188
rect 25004 54176 25010 54188
rect 25041 54179 25099 54185
rect 25041 54176 25053 54179
rect 25004 54148 25053 54176
rect 25004 54136 25010 54148
rect 25041 54145 25053 54148
rect 25087 54145 25099 54179
rect 26326 54176 26332 54188
rect 26287 54148 26332 54176
rect 25041 54139 25099 54145
rect 26326 54136 26332 54148
rect 26384 54136 26390 54188
rect 27062 54136 27068 54188
rect 27120 54176 27126 54188
rect 27229 54179 27287 54185
rect 27229 54176 27241 54179
rect 27120 54148 27241 54176
rect 27120 54136 27126 54148
rect 27229 54145 27241 54148
rect 27275 54145 27287 54179
rect 29822 54176 29828 54188
rect 29783 54148 29828 54176
rect 27229 54139 27287 54145
rect 29822 54136 29828 54148
rect 29880 54136 29886 54188
rect 30092 54179 30150 54185
rect 30092 54145 30104 54179
rect 30138 54176 30150 54179
rect 30650 54176 30656 54188
rect 30138 54148 30656 54176
rect 30138 54145 30150 54148
rect 30092 54139 30150 54145
rect 30650 54136 30656 54148
rect 30708 54136 30714 54188
rect 20680 54080 22324 54108
rect 26421 54111 26479 54117
rect 20680 54068 20686 54080
rect 26421 54077 26433 54111
rect 26467 54108 26479 54111
rect 26973 54111 27031 54117
rect 26973 54108 26985 54111
rect 26467 54080 26985 54108
rect 26467 54077 26479 54080
rect 26421 54071 26479 54077
rect 26973 54077 26985 54080
rect 27019 54077 27031 54111
rect 31726 54108 31754 54216
rect 37820 54213 37832 54247
rect 37866 54244 37878 54247
rect 38286 54244 38292 54256
rect 37866 54216 38292 54244
rect 37866 54213 37878 54216
rect 37820 54207 37878 54213
rect 38286 54204 38292 54216
rect 38344 54204 38350 54256
rect 41386 54244 41414 54284
rect 45186 54272 45192 54284
rect 45244 54272 45250 54324
rect 45646 54312 45652 54324
rect 45607 54284 45652 54312
rect 45646 54272 45652 54284
rect 45704 54272 45710 54324
rect 47670 54272 47676 54324
rect 47728 54312 47734 54324
rect 47765 54315 47823 54321
rect 47765 54312 47777 54315
rect 47728 54284 47777 54312
rect 47728 54272 47734 54284
rect 47765 54281 47777 54284
rect 47811 54281 47823 54315
rect 47765 54275 47823 54281
rect 48498 54272 48504 54324
rect 48556 54312 48562 54324
rect 48961 54315 49019 54321
rect 48961 54312 48973 54315
rect 48556 54284 48973 54312
rect 48556 54272 48562 54284
rect 48961 54281 48973 54284
rect 49007 54281 49019 54315
rect 48961 54275 49019 54281
rect 50249 54315 50307 54321
rect 50249 54281 50261 54315
rect 50295 54312 50307 54315
rect 51258 54312 51264 54324
rect 50295 54284 51264 54312
rect 50295 54281 50307 54284
rect 50249 54275 50307 54281
rect 51258 54272 51264 54284
rect 51316 54272 51322 54324
rect 40144 54216 41414 54244
rect 43456 54216 45876 54244
rect 32392 54179 32450 54185
rect 32392 54145 32404 54179
rect 32438 54176 32450 54179
rect 32858 54176 32864 54188
rect 32438 54148 32864 54176
rect 32438 54145 32450 54148
rect 32392 54139 32450 54145
rect 32858 54136 32864 54148
rect 32916 54136 32922 54188
rect 37550 54176 37556 54188
rect 37511 54148 37556 54176
rect 37550 54136 37556 54148
rect 37608 54136 37614 54188
rect 40034 54176 40040 54188
rect 39995 54148 40040 54176
rect 40034 54136 40040 54148
rect 40092 54136 40098 54188
rect 40144 54185 40172 54216
rect 40129 54179 40187 54185
rect 40129 54145 40141 54179
rect 40175 54145 40187 54179
rect 40129 54139 40187 54145
rect 40313 54179 40371 54185
rect 40313 54145 40325 54179
rect 40359 54176 40371 54179
rect 40957 54179 41015 54185
rect 40957 54176 40969 54179
rect 40359 54148 40969 54176
rect 40359 54145 40371 54148
rect 40313 54139 40371 54145
rect 40957 54145 40969 54148
rect 41003 54145 41015 54179
rect 40957 54139 41015 54145
rect 32125 54111 32183 54117
rect 32125 54108 32137 54111
rect 31726 54080 32137 54108
rect 26973 54071 27031 54077
rect 32125 54077 32137 54080
rect 32171 54077 32183 54111
rect 40144 54108 40172 54139
rect 41414 54136 41420 54188
rect 41472 54176 41478 54188
rect 41472 54148 41517 54176
rect 41472 54136 41478 54148
rect 32125 54071 32183 54077
rect 38764 54080 40172 54108
rect 17954 54040 17960 54052
rect 17915 54012 17960 54040
rect 17954 54000 17960 54012
rect 18012 54000 18018 54052
rect 24581 54043 24639 54049
rect 24581 54009 24593 54043
rect 24627 54040 24639 54043
rect 29178 54040 29184 54052
rect 24627 54012 25636 54040
rect 24627 54009 24639 54012
rect 24581 54003 24639 54009
rect 1946 53972 1952 53984
rect 1907 53944 1952 53972
rect 1946 53932 1952 53944
rect 2004 53932 2010 53984
rect 16117 53975 16175 53981
rect 16117 53941 16129 53975
rect 16163 53972 16175 53975
rect 16850 53972 16856 53984
rect 16163 53944 16856 53972
rect 16163 53941 16175 53944
rect 16117 53935 16175 53941
rect 16850 53932 16856 53944
rect 16908 53932 16914 53984
rect 16942 53932 16948 53984
rect 17000 53972 17006 53984
rect 18322 53972 18328 53984
rect 17000 53944 18328 53972
rect 17000 53932 17006 53944
rect 18322 53932 18328 53944
rect 18380 53932 18386 53984
rect 19334 53932 19340 53984
rect 19392 53972 19398 53984
rect 20993 53975 21051 53981
rect 20993 53972 21005 53975
rect 19392 53944 21005 53972
rect 19392 53932 19398 53944
rect 20993 53941 21005 53944
rect 21039 53941 21051 53975
rect 20993 53935 21051 53941
rect 22830 53932 22836 53984
rect 22888 53972 22894 53984
rect 24596 53972 24624 54003
rect 22888 53944 24624 53972
rect 22888 53932 22894 53944
rect 24854 53932 24860 53984
rect 24912 53972 24918 53984
rect 25041 53975 25099 53981
rect 25041 53972 25053 53975
rect 24912 53944 25053 53972
rect 24912 53932 24918 53944
rect 25041 53941 25053 53944
rect 25087 53941 25099 53975
rect 25608 53972 25636 54012
rect 27908 54012 29184 54040
rect 27908 53972 27936 54012
rect 29178 54000 29184 54012
rect 29236 54000 29242 54052
rect 28350 53972 28356 53984
rect 25608 53944 27936 53972
rect 28311 53944 28356 53972
rect 25041 53935 25099 53941
rect 28350 53932 28356 53944
rect 28408 53932 28414 53984
rect 29822 53932 29828 53984
rect 29880 53972 29886 53984
rect 31205 53975 31263 53981
rect 31205 53972 31217 53975
rect 29880 53944 31217 53972
rect 29880 53932 29886 53944
rect 31205 53941 31217 53944
rect 31251 53941 31263 53975
rect 32140 53972 32168 54071
rect 32766 53972 32772 53984
rect 32140 53944 32772 53972
rect 31205 53935 31263 53941
rect 32766 53932 32772 53944
rect 32824 53932 32830 53984
rect 37826 53932 37832 53984
rect 37884 53972 37890 53984
rect 38764 53972 38792 54080
rect 41322 54000 41328 54052
rect 41380 54040 41386 54052
rect 43456 54040 43484 54216
rect 43622 54176 43628 54188
rect 43583 54148 43628 54176
rect 43622 54136 43628 54148
rect 43680 54136 43686 54188
rect 43714 54136 43720 54188
rect 43772 54176 43778 54188
rect 45848 54185 45876 54216
rect 43881 54179 43939 54185
rect 43881 54176 43893 54179
rect 43772 54148 43893 54176
rect 43772 54136 43778 54148
rect 43881 54145 43893 54148
rect 43927 54145 43939 54179
rect 43881 54139 43939 54145
rect 45833 54179 45891 54185
rect 45833 54145 45845 54179
rect 45879 54145 45891 54179
rect 45833 54139 45891 54145
rect 46934 54136 46940 54188
rect 46992 54176 46998 54188
rect 47581 54179 47639 54185
rect 47581 54176 47593 54179
rect 46992 54148 47593 54176
rect 46992 54136 46998 54148
rect 47581 54145 47593 54148
rect 47627 54145 47639 54179
rect 48682 54176 48688 54188
rect 48643 54148 48688 54176
rect 47581 54139 47639 54145
rect 48682 54136 48688 54148
rect 48740 54136 48746 54188
rect 48777 54179 48835 54185
rect 48777 54145 48789 54179
rect 48823 54176 48835 54179
rect 49694 54176 49700 54188
rect 48823 54148 49700 54176
rect 48823 54145 48835 54148
rect 48777 54139 48835 54145
rect 49694 54136 49700 54148
rect 49752 54176 49758 54188
rect 50062 54176 50068 54188
rect 49752 54148 50068 54176
rect 49752 54136 49758 54148
rect 50062 54136 50068 54148
rect 50120 54136 50126 54188
rect 50154 54136 50160 54188
rect 50212 54176 50218 54188
rect 50893 54179 50951 54185
rect 50893 54176 50905 54179
rect 50212 54148 50905 54176
rect 50212 54136 50218 54148
rect 50893 54145 50905 54148
rect 50939 54145 50951 54179
rect 50893 54139 50951 54145
rect 46109 54111 46167 54117
rect 46109 54077 46121 54111
rect 46155 54108 46167 54111
rect 46566 54108 46572 54120
rect 46155 54080 46572 54108
rect 46155 54077 46167 54080
rect 46109 54071 46167 54077
rect 46566 54068 46572 54080
rect 46624 54068 46630 54120
rect 49878 54108 49884 54120
rect 49839 54080 49884 54108
rect 49878 54068 49884 54080
rect 49936 54068 49942 54120
rect 41380 54012 43484 54040
rect 41380 54000 41386 54012
rect 38930 53972 38936 53984
rect 37884 53944 38792 53972
rect 38891 53944 38936 53972
rect 37884 53932 37890 53944
rect 38930 53932 38936 53944
rect 38988 53932 38994 53984
rect 40770 53972 40776 53984
rect 40731 53944 40776 53972
rect 40770 53932 40776 53944
rect 40828 53932 40834 53984
rect 41506 53972 41512 53984
rect 41467 53944 41512 53972
rect 41506 53932 41512 53944
rect 41564 53932 41570 53984
rect 45005 53975 45063 53981
rect 45005 53941 45017 53975
rect 45051 53972 45063 53975
rect 45462 53972 45468 53984
rect 45051 53944 45468 53972
rect 45051 53941 45063 53944
rect 45005 53935 45063 53941
rect 45462 53932 45468 53944
rect 45520 53932 45526 53984
rect 45554 53932 45560 53984
rect 45612 53972 45618 53984
rect 46017 53975 46075 53981
rect 46017 53972 46029 53975
rect 45612 53944 46029 53972
rect 45612 53932 45618 53944
rect 46017 53941 46029 53944
rect 46063 53941 46075 53975
rect 46017 53935 46075 53941
rect 50709 53975 50767 53981
rect 50709 53941 50721 53975
rect 50755 53972 50767 53975
rect 50798 53972 50804 53984
rect 50755 53944 50804 53972
rect 50755 53941 50767 53944
rect 50709 53935 50767 53941
rect 50798 53932 50804 53944
rect 50856 53932 50862 53984
rect 1104 53882 68816 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 65654 53882
rect 65706 53830 65718 53882
rect 65770 53830 65782 53882
rect 65834 53830 65846 53882
rect 65898 53830 65910 53882
rect 65962 53830 68816 53882
rect 1104 53808 68816 53830
rect 6089 53771 6147 53777
rect 6089 53737 6101 53771
rect 6135 53768 6147 53771
rect 6546 53768 6552 53780
rect 6135 53740 6552 53768
rect 6135 53737 6147 53740
rect 6089 53731 6147 53737
rect 6546 53728 6552 53740
rect 6604 53728 6610 53780
rect 16942 53768 16948 53780
rect 16903 53740 16948 53768
rect 16942 53728 16948 53740
rect 17000 53728 17006 53780
rect 19981 53771 20039 53777
rect 19981 53737 19993 53771
rect 20027 53737 20039 53771
rect 19981 53731 20039 53737
rect 20165 53771 20223 53777
rect 20165 53737 20177 53771
rect 20211 53768 20223 53771
rect 20346 53768 20352 53780
rect 20211 53740 20352 53768
rect 20211 53737 20223 53740
rect 20165 53731 20223 53737
rect 19996 53700 20024 53731
rect 20346 53728 20352 53740
rect 20404 53728 20410 53780
rect 21545 53771 21603 53777
rect 21545 53737 21557 53771
rect 21591 53768 21603 53771
rect 23382 53768 23388 53780
rect 21591 53740 23388 53768
rect 21591 53737 21603 53740
rect 21545 53731 21603 53737
rect 23382 53728 23388 53740
rect 23440 53728 23446 53780
rect 26973 53771 27031 53777
rect 26973 53737 26985 53771
rect 27019 53768 27031 53771
rect 27062 53768 27068 53780
rect 27019 53740 27068 53768
rect 27019 53737 27031 53740
rect 26973 53731 27031 53737
rect 27062 53728 27068 53740
rect 27120 53728 27126 53780
rect 27246 53728 27252 53780
rect 27304 53768 27310 53780
rect 30006 53768 30012 53780
rect 27304 53740 29868 53768
rect 29919 53740 30012 53768
rect 27304 53728 27310 53740
rect 20438 53700 20444 53712
rect 19996 53672 20444 53700
rect 20438 53660 20444 53672
rect 20496 53660 20502 53712
rect 26234 53700 26240 53712
rect 26147 53672 26240 53700
rect 26234 53660 26240 53672
rect 26292 53700 26298 53712
rect 29086 53700 29092 53712
rect 26292 53672 29092 53700
rect 26292 53660 26298 53672
rect 29086 53660 29092 53672
rect 29144 53660 29150 53712
rect 1397 53635 1455 53641
rect 1397 53601 1409 53635
rect 1443 53632 1455 53635
rect 1946 53632 1952 53644
rect 1443 53604 1952 53632
rect 1443 53601 1455 53604
rect 1397 53595 1455 53601
rect 1946 53592 1952 53604
rect 2004 53592 2010 53644
rect 2774 53632 2780 53644
rect 2735 53604 2780 53632
rect 2774 53592 2780 53604
rect 2832 53592 2838 53644
rect 15194 53632 15200 53644
rect 14660 53604 15200 53632
rect 5997 53567 6055 53573
rect 5997 53533 6009 53567
rect 6043 53564 6055 53567
rect 6362 53564 6368 53576
rect 6043 53536 6368 53564
rect 6043 53533 6055 53536
rect 5997 53527 6055 53533
rect 6362 53524 6368 53536
rect 6420 53524 6426 53576
rect 13449 53567 13507 53573
rect 13449 53533 13461 53567
rect 13495 53564 13507 53567
rect 13814 53564 13820 53576
rect 13495 53536 13820 53564
rect 13495 53533 13507 53536
rect 13449 53527 13507 53533
rect 13814 53524 13820 53536
rect 13872 53524 13878 53576
rect 14660 53573 14688 53604
rect 15194 53592 15200 53604
rect 15252 53592 15258 53644
rect 22186 53592 22192 53644
rect 22244 53632 22250 53644
rect 22741 53635 22799 53641
rect 22741 53632 22753 53635
rect 22244 53604 22753 53632
rect 22244 53592 22250 53604
rect 22741 53601 22753 53604
rect 22787 53601 22799 53635
rect 24854 53632 24860 53644
rect 24815 53604 24860 53632
rect 22741 53595 22799 53601
rect 24854 53592 24860 53604
rect 24912 53592 24918 53644
rect 27985 53635 28043 53641
rect 27985 53632 27997 53635
rect 27172 53604 27997 53632
rect 14553 53567 14611 53573
rect 14553 53533 14565 53567
rect 14599 53533 14611 53567
rect 14553 53527 14611 53533
rect 14645 53567 14703 53573
rect 14645 53533 14657 53567
rect 14691 53533 14703 53567
rect 15562 53564 15568 53576
rect 15523 53536 15568 53564
rect 14645 53527 14703 53533
rect 1581 53499 1639 53505
rect 1581 53465 1593 53499
rect 1627 53496 1639 53499
rect 2406 53496 2412 53508
rect 1627 53468 2412 53496
rect 1627 53465 1639 53468
rect 1581 53459 1639 53465
rect 2406 53456 2412 53468
rect 2464 53456 2470 53508
rect 14568 53496 14596 53527
rect 15562 53524 15568 53536
rect 15620 53524 15626 53576
rect 17402 53564 17408 53576
rect 17363 53536 17408 53564
rect 17402 53524 17408 53536
rect 17460 53524 17466 53576
rect 21726 53564 21732 53576
rect 20027 53533 20085 53539
rect 21687 53536 21732 53564
rect 15194 53496 15200 53508
rect 14568 53468 15200 53496
rect 15194 53456 15200 53468
rect 15252 53456 15258 53508
rect 15832 53499 15890 53505
rect 15832 53465 15844 53499
rect 15878 53496 15890 53499
rect 16666 53496 16672 53508
rect 15878 53468 16672 53496
rect 15878 53465 15890 53468
rect 15832 53459 15890 53465
rect 16666 53456 16672 53468
rect 16724 53456 16730 53508
rect 18509 53499 18567 53505
rect 18509 53465 18521 53499
rect 18555 53496 18567 53499
rect 18874 53496 18880 53508
rect 18555 53468 18880 53496
rect 18555 53465 18567 53468
rect 18509 53459 18567 53465
rect 18874 53456 18880 53468
rect 18932 53456 18938 53508
rect 19334 53456 19340 53508
rect 19392 53496 19398 53508
rect 19797 53499 19855 53505
rect 19797 53496 19809 53499
rect 19392 53468 19809 53496
rect 19392 53456 19398 53468
rect 19797 53465 19809 53468
rect 19843 53465 19855 53499
rect 20027 53499 20039 53533
rect 20073 53530 20085 53533
rect 20073 53508 20107 53530
rect 21726 53524 21732 53536
rect 21784 53524 21790 53576
rect 25130 53573 25136 53576
rect 22005 53567 22063 53573
rect 22005 53564 22017 53567
rect 21836 53536 22017 53564
rect 20073 53499 20076 53508
rect 20027 53493 20076 53499
rect 19797 53459 19855 53465
rect 20070 53456 20076 53493
rect 20128 53456 20134 53508
rect 20162 53456 20168 53508
rect 20220 53496 20226 53508
rect 21836 53496 21864 53536
rect 22005 53533 22017 53536
rect 22051 53533 22063 53567
rect 22005 53527 22063 53533
rect 22465 53567 22523 53573
rect 22465 53533 22477 53567
rect 22511 53533 22523 53567
rect 25124 53564 25136 53573
rect 25091 53536 25136 53564
rect 22465 53527 22523 53533
rect 25124 53527 25136 53536
rect 20220 53468 21864 53496
rect 21913 53499 21971 53505
rect 20220 53456 20226 53468
rect 21913 53465 21925 53499
rect 21959 53496 21971 53499
rect 22186 53496 22192 53508
rect 21959 53468 22192 53496
rect 21959 53465 21971 53468
rect 21913 53459 21971 53465
rect 22186 53456 22192 53468
rect 22244 53456 22250 53508
rect 13449 53431 13507 53437
rect 13449 53397 13461 53431
rect 13495 53428 13507 53431
rect 13538 53428 13544 53440
rect 13495 53400 13544 53428
rect 13495 53397 13507 53400
rect 13449 53391 13507 53397
rect 13538 53388 13544 53400
rect 13596 53388 13602 53440
rect 14274 53388 14280 53440
rect 14332 53428 14338 53440
rect 14829 53431 14887 53437
rect 14829 53428 14841 53431
rect 14332 53400 14841 53428
rect 14332 53388 14338 53400
rect 14829 53397 14841 53400
rect 14875 53397 14887 53431
rect 14829 53391 14887 53397
rect 17310 53388 17316 53440
rect 17368 53428 17374 53440
rect 17589 53431 17647 53437
rect 17589 53428 17601 53431
rect 17368 53400 17601 53428
rect 17368 53388 17374 53400
rect 17589 53397 17601 53400
rect 17635 53397 17647 53431
rect 18598 53428 18604 53440
rect 18559 53400 18604 53428
rect 17589 53391 17647 53397
rect 18598 53388 18604 53400
rect 18656 53388 18662 53440
rect 22480 53428 22508 53527
rect 25130 53524 25136 53527
rect 25188 53524 25194 53576
rect 27172 53573 27200 53604
rect 27985 53601 27997 53604
rect 28031 53601 28043 53635
rect 29840 53632 29868 53740
rect 30006 53728 30012 53740
rect 30064 53768 30070 53780
rect 30282 53768 30288 53780
rect 30064 53740 30288 53768
rect 30064 53728 30070 53740
rect 30282 53728 30288 53740
rect 30340 53728 30346 53780
rect 30650 53768 30656 53780
rect 30611 53740 30656 53768
rect 30650 53728 30656 53740
rect 30708 53728 30714 53780
rect 32858 53768 32864 53780
rect 32819 53740 32864 53768
rect 32858 53728 32864 53740
rect 32916 53728 32922 53780
rect 37458 53728 37464 53780
rect 37516 53768 37522 53780
rect 43530 53768 43536 53780
rect 37516 53740 43536 53768
rect 37516 53728 37522 53740
rect 43530 53728 43536 53740
rect 43588 53728 43594 53780
rect 43625 53771 43683 53777
rect 43625 53737 43637 53771
rect 43671 53768 43683 53771
rect 43714 53768 43720 53780
rect 43671 53740 43720 53768
rect 43671 53737 43683 53740
rect 43625 53731 43683 53737
rect 43714 53728 43720 53740
rect 43772 53728 43778 53780
rect 45281 53771 45339 53777
rect 45281 53737 45293 53771
rect 45327 53768 45339 53771
rect 45830 53768 45836 53780
rect 45327 53740 45836 53768
rect 45327 53737 45339 53740
rect 45281 53731 45339 53737
rect 45830 53728 45836 53740
rect 45888 53768 45894 53780
rect 47578 53768 47584 53780
rect 45888 53740 47584 53768
rect 45888 53728 45894 53740
rect 47578 53728 47584 53740
rect 47636 53728 47642 53780
rect 48682 53768 48688 53780
rect 48643 53740 48688 53768
rect 48682 53728 48688 53740
rect 48740 53728 48746 53780
rect 30098 53660 30104 53712
rect 30156 53700 30162 53712
rect 48593 53703 48651 53709
rect 30156 53672 36124 53700
rect 30156 53660 30162 53672
rect 31588 53641 31616 53672
rect 31573 53635 31631 53641
rect 29840 53604 30972 53632
rect 27985 53595 28043 53601
rect 27157 53567 27215 53573
rect 27157 53533 27169 53567
rect 27203 53533 27215 53567
rect 27157 53527 27215 53533
rect 27709 53567 27767 53573
rect 27709 53533 27721 53567
rect 27755 53533 27767 53567
rect 27709 53527 27767 53533
rect 22554 53456 22560 53508
rect 22612 53496 22618 53508
rect 27246 53496 27252 53508
rect 22612 53468 27252 53496
rect 22612 53456 22618 53468
rect 27246 53456 27252 53468
rect 27304 53456 27310 53508
rect 27724 53496 27752 53527
rect 27798 53524 27804 53576
rect 27856 53564 27862 53576
rect 27856 53536 27901 53564
rect 27856 53524 27862 53536
rect 29730 53524 29736 53576
rect 29788 53564 29794 53576
rect 30837 53567 30895 53573
rect 29788 53539 30098 53564
rect 29788 53536 30113 53539
rect 29788 53524 29794 53536
rect 30055 53533 30113 53536
rect 28350 53496 28356 53508
rect 27724 53468 28356 53496
rect 28350 53456 28356 53468
rect 28408 53456 28414 53508
rect 29822 53496 29828 53508
rect 29783 53468 29828 53496
rect 29822 53456 29828 53468
rect 29880 53456 29886 53508
rect 30055 53499 30067 53533
rect 30101 53499 30113 53533
rect 30837 53533 30849 53567
rect 30883 53533 30895 53567
rect 30944 53564 30972 53604
rect 31573 53601 31585 53635
rect 31619 53601 31631 53635
rect 31573 53595 31631 53601
rect 31754 53592 31760 53644
rect 31812 53632 31818 53644
rect 31849 53635 31907 53641
rect 31849 53632 31861 53635
rect 31812 53604 31861 53632
rect 31812 53592 31818 53604
rect 31849 53601 31861 53604
rect 31895 53601 31907 53635
rect 31849 53595 31907 53601
rect 35069 53635 35127 53641
rect 35069 53601 35081 53635
rect 35115 53632 35127 53635
rect 35434 53632 35440 53644
rect 35115 53604 35440 53632
rect 35115 53601 35127 53604
rect 35069 53595 35127 53601
rect 35434 53592 35440 53604
rect 35492 53592 35498 53644
rect 32398 53564 32404 53576
rect 30944 53536 32404 53564
rect 30837 53527 30895 53533
rect 30055 53493 30113 53499
rect 30098 53428 30104 53440
rect 22480 53400 30104 53428
rect 30098 53388 30104 53400
rect 30156 53388 30162 53440
rect 30193 53431 30251 53437
rect 30193 53397 30205 53431
rect 30239 53428 30251 53431
rect 30852 53428 30880 53527
rect 32398 53524 32404 53536
rect 32456 53524 32462 53576
rect 33134 53564 33140 53576
rect 33095 53536 33140 53564
rect 33134 53524 33140 53536
rect 33192 53524 33198 53576
rect 33229 53567 33287 53573
rect 33229 53533 33241 53567
rect 33275 53533 33287 53567
rect 33229 53527 33287 53533
rect 33244 53496 33272 53527
rect 33318 53524 33324 53576
rect 33376 53564 33382 53576
rect 33505 53567 33563 53573
rect 33376 53536 33421 53564
rect 33376 53524 33382 53536
rect 33505 53533 33517 53567
rect 33551 53564 33563 53567
rect 35250 53564 35256 53576
rect 33551 53536 34652 53564
rect 35211 53536 35256 53564
rect 33551 53533 33563 53536
rect 33505 53527 33563 53533
rect 34422 53496 34428 53508
rect 33244 53468 34428 53496
rect 34422 53456 34428 53468
rect 34480 53456 34486 53508
rect 30239 53400 30880 53428
rect 34624 53428 34652 53536
rect 35250 53524 35256 53536
rect 35308 53524 35314 53576
rect 35529 53567 35587 53573
rect 35529 53533 35541 53567
rect 35575 53564 35587 53567
rect 35618 53564 35624 53576
rect 35575 53536 35624 53564
rect 35575 53533 35587 53536
rect 35529 53527 35587 53533
rect 35618 53524 35624 53536
rect 35676 53564 35682 53576
rect 35986 53564 35992 53576
rect 35676 53536 35992 53564
rect 35676 53524 35682 53536
rect 35986 53524 35992 53536
rect 36044 53524 36050 53576
rect 35437 53499 35495 53505
rect 35437 53465 35449 53499
rect 35483 53496 35495 53499
rect 35710 53496 35716 53508
rect 35483 53468 35716 53496
rect 35483 53465 35495 53468
rect 35437 53459 35495 53465
rect 35710 53456 35716 53468
rect 35768 53456 35774 53508
rect 35894 53428 35900 53440
rect 34624 53400 35900 53428
rect 30239 53397 30251 53400
rect 30193 53391 30251 53397
rect 35894 53388 35900 53400
rect 35952 53388 35958 53440
rect 36096 53428 36124 53672
rect 48593 53669 48605 53703
rect 48639 53700 48651 53703
rect 49878 53700 49884 53712
rect 48639 53672 49884 53700
rect 48639 53669 48651 53672
rect 48593 53663 48651 53669
rect 49878 53660 49884 53672
rect 49936 53660 49942 53712
rect 41506 53632 41512 53644
rect 41467 53604 41512 53632
rect 41506 53592 41512 53604
rect 41564 53592 41570 53644
rect 43162 53592 43168 53644
rect 43220 53632 43226 53644
rect 45186 53632 45192 53644
rect 43220 53604 45192 53632
rect 43220 53592 43226 53604
rect 36541 53567 36599 53573
rect 36541 53533 36553 53567
rect 36587 53564 36599 53567
rect 37550 53564 37556 53576
rect 36587 53536 37556 53564
rect 36587 53533 36599 53536
rect 36541 53527 36599 53533
rect 37550 53524 37556 53536
rect 37608 53524 37614 53576
rect 39209 53567 39267 53573
rect 39209 53533 39221 53567
rect 39255 53564 39267 53567
rect 39390 53564 39396 53576
rect 39255 53536 39396 53564
rect 39255 53533 39267 53536
rect 39209 53527 39267 53533
rect 39390 53524 39396 53536
rect 39448 53564 39454 53576
rect 40681 53567 40739 53573
rect 40681 53564 40693 53567
rect 39448 53536 40693 53564
rect 39448 53524 39454 53536
rect 40681 53533 40693 53536
rect 40727 53564 40739 53567
rect 41414 53564 41420 53576
rect 40727 53536 41420 53564
rect 40727 53533 40739 53536
rect 40681 53527 40739 53533
rect 41414 53524 41420 53536
rect 41472 53524 41478 53576
rect 43625 53567 43683 53573
rect 43625 53533 43637 53567
rect 43671 53564 43683 53567
rect 43714 53564 43720 53576
rect 43671 53536 43720 53564
rect 43671 53533 43683 53536
rect 43625 53527 43683 53533
rect 43714 53524 43720 53536
rect 43772 53524 43778 53576
rect 43824 53573 43852 53604
rect 45186 53592 45192 53604
rect 45244 53592 45250 53644
rect 46566 53592 46572 53644
rect 46624 53632 46630 53644
rect 46624 53604 48820 53632
rect 46624 53592 46630 53604
rect 43809 53567 43867 53573
rect 43809 53533 43821 53567
rect 43855 53533 43867 53567
rect 43809 53527 43867 53533
rect 45097 53567 45155 53573
rect 45097 53533 45109 53567
rect 45143 53533 45155 53567
rect 45097 53527 45155 53533
rect 36808 53499 36866 53505
rect 36808 53465 36820 53499
rect 36854 53496 36866 53499
rect 37274 53496 37280 53508
rect 36854 53468 37280 53496
rect 36854 53465 36866 53468
rect 36808 53459 36866 53465
rect 37274 53456 37280 53468
rect 37332 53456 37338 53508
rect 38838 53496 38844 53508
rect 37384 53468 38844 53496
rect 37384 53428 37412 53468
rect 38838 53456 38844 53468
rect 38896 53456 38902 53508
rect 40218 53456 40224 53508
rect 40276 53496 40282 53508
rect 41782 53505 41788 53508
rect 40313 53499 40371 53505
rect 40313 53496 40325 53499
rect 40276 53468 40325 53496
rect 40276 53456 40282 53468
rect 40313 53465 40325 53468
rect 40359 53496 40371 53499
rect 40359 53468 41414 53496
rect 40359 53465 40371 53468
rect 40313 53459 40371 53465
rect 37918 53428 37924 53440
rect 36096 53400 37412 53428
rect 37879 53400 37924 53428
rect 37918 53388 37924 53400
rect 37976 53388 37982 53440
rect 39209 53431 39267 53437
rect 39209 53397 39221 53431
rect 39255 53428 39267 53431
rect 39482 53428 39488 53440
rect 39255 53400 39488 53428
rect 39255 53397 39267 53400
rect 39209 53391 39267 53397
rect 39482 53388 39488 53400
rect 39540 53388 39546 53440
rect 41386 53428 41414 53468
rect 41776 53459 41788 53505
rect 41840 53496 41846 53508
rect 45002 53496 45008 53508
rect 41840 53468 41876 53496
rect 42720 53468 45008 53496
rect 41782 53456 41788 53459
rect 41840 53456 41846 53468
rect 42720 53428 42748 53468
rect 45002 53456 45008 53468
rect 45060 53496 45066 53508
rect 45112 53496 45140 53527
rect 46106 53524 46112 53576
rect 46164 53564 46170 53576
rect 46201 53567 46259 53573
rect 46201 53564 46213 53567
rect 46164 53536 46213 53564
rect 46164 53524 46170 53536
rect 46201 53533 46213 53536
rect 46247 53533 46259 53567
rect 46201 53527 46259 53533
rect 46385 53567 46443 53573
rect 46385 53533 46397 53567
rect 46431 53533 46443 53567
rect 48498 53564 48504 53576
rect 48459 53536 48504 53564
rect 46385 53527 46443 53533
rect 46400 53496 46428 53527
rect 48498 53524 48504 53536
rect 48556 53524 48562 53576
rect 48792 53573 48820 53604
rect 48777 53567 48835 53573
rect 48777 53533 48789 53567
rect 48823 53533 48835 53567
rect 48777 53527 48835 53533
rect 50525 53567 50583 53573
rect 50525 53533 50537 53567
rect 50571 53564 50583 53567
rect 50614 53564 50620 53576
rect 50571 53536 50620 53564
rect 50571 53533 50583 53536
rect 50525 53527 50583 53533
rect 50614 53524 50620 53536
rect 50672 53524 50678 53576
rect 50798 53573 50804 53576
rect 50792 53564 50804 53573
rect 50759 53536 50804 53564
rect 50792 53527 50804 53536
rect 50798 53524 50804 53527
rect 50856 53524 50862 53576
rect 45060 53468 45140 53496
rect 46216 53468 46428 53496
rect 45060 53456 45066 53468
rect 46216 53440 46244 53468
rect 48222 53456 48228 53508
rect 48280 53496 48286 53508
rect 48317 53499 48375 53505
rect 48317 53496 48329 53499
rect 48280 53468 48329 53496
rect 48280 53456 48286 53468
rect 48317 53465 48329 53468
rect 48363 53465 48375 53499
rect 48317 53459 48375 53465
rect 42886 53428 42892 53440
rect 41386 53400 42748 53428
rect 42847 53400 42892 53428
rect 42886 53388 42892 53400
rect 42944 53388 42950 53440
rect 46198 53388 46204 53440
rect 46256 53388 46262 53440
rect 46382 53428 46388 53440
rect 46343 53400 46388 53428
rect 46382 53388 46388 53400
rect 46440 53388 46446 53440
rect 48869 53431 48927 53437
rect 48869 53397 48881 53431
rect 48915 53428 48927 53431
rect 48958 53428 48964 53440
rect 48915 53400 48964 53428
rect 48915 53397 48927 53400
rect 48869 53391 48927 53397
rect 48958 53388 48964 53400
rect 49016 53388 49022 53440
rect 49878 53388 49884 53440
rect 49936 53428 49942 53440
rect 51905 53431 51963 53437
rect 51905 53428 51917 53431
rect 49936 53400 51917 53428
rect 49936 53388 49942 53400
rect 51905 53397 51917 53400
rect 51951 53397 51963 53431
rect 51905 53391 51963 53397
rect 1104 53338 68816 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 68816 53338
rect 1104 53264 68816 53286
rect 2406 53224 2412 53236
rect 2367 53196 2412 53224
rect 2406 53184 2412 53196
rect 2464 53184 2470 53236
rect 15562 53184 15568 53236
rect 15620 53224 15626 53236
rect 15749 53227 15807 53233
rect 15749 53224 15761 53227
rect 15620 53196 15761 53224
rect 15620 53184 15626 53196
rect 15749 53193 15761 53196
rect 15795 53193 15807 53227
rect 16666 53224 16672 53236
rect 16627 53196 16672 53224
rect 15749 53187 15807 53193
rect 16666 53184 16672 53196
rect 16724 53184 16730 53236
rect 17402 53184 17408 53236
rect 17460 53224 17466 53236
rect 22922 53224 22928 53236
rect 17460 53196 22928 53224
rect 17460 53184 17466 53196
rect 22922 53184 22928 53196
rect 22980 53224 22986 53236
rect 23290 53224 23296 53236
rect 22980 53196 23296 53224
rect 22980 53184 22986 53196
rect 23290 53184 23296 53196
rect 23348 53184 23354 53236
rect 25406 53184 25412 53236
rect 25464 53224 25470 53236
rect 25685 53227 25743 53233
rect 25685 53224 25697 53227
rect 25464 53196 25697 53224
rect 25464 53184 25470 53196
rect 25685 53193 25697 53196
rect 25731 53193 25743 53227
rect 29917 53227 29975 53233
rect 25685 53187 25743 53193
rect 26436 53196 29776 53224
rect 16758 53116 16764 53168
rect 16816 53156 16822 53168
rect 24854 53156 24860 53168
rect 16816 53128 24860 53156
rect 16816 53116 16822 53128
rect 24854 53116 24860 53128
rect 24912 53116 24918 53168
rect 26234 53156 26240 53168
rect 25424 53128 26240 53156
rect 2317 53091 2375 53097
rect 2317 53057 2329 53091
rect 2363 53088 2375 53091
rect 5166 53088 5172 53100
rect 2363 53060 5172 53088
rect 2363 53057 2375 53060
rect 2317 53051 2375 53057
rect 5166 53048 5172 53060
rect 5224 53048 5230 53100
rect 13538 53088 13544 53100
rect 13499 53060 13544 53088
rect 13538 53048 13544 53060
rect 13596 53048 13602 53100
rect 13808 53091 13866 53097
rect 13808 53057 13820 53091
rect 13854 53088 13866 53091
rect 14090 53088 14096 53100
rect 13854 53060 14096 53088
rect 13854 53057 13866 53060
rect 13808 53051 13866 53057
rect 14090 53048 14096 53060
rect 14148 53048 14154 53100
rect 15749 53091 15807 53097
rect 15749 53057 15761 53091
rect 15795 53088 15807 53091
rect 15838 53088 15844 53100
rect 15795 53060 15844 53088
rect 15795 53057 15807 53060
rect 15749 53051 15807 53057
rect 15838 53048 15844 53060
rect 15896 53048 15902 53100
rect 16850 53088 16856 53100
rect 16811 53060 16856 53088
rect 16850 53048 16856 53060
rect 16908 53048 16914 53100
rect 19521 53091 19579 53097
rect 19521 53057 19533 53091
rect 19567 53088 19579 53091
rect 19978 53088 19984 53100
rect 19567 53060 19984 53088
rect 19567 53057 19579 53060
rect 19521 53051 19579 53057
rect 19978 53048 19984 53060
rect 20036 53048 20042 53100
rect 20809 53091 20867 53097
rect 20809 53057 20821 53091
rect 20855 53088 20867 53091
rect 20898 53088 20904 53100
rect 20855 53060 20904 53088
rect 20855 53057 20867 53060
rect 20809 53051 20867 53057
rect 20898 53048 20904 53060
rect 20956 53048 20962 53100
rect 21726 53048 21732 53100
rect 21784 53088 21790 53100
rect 22649 53091 22707 53097
rect 22649 53088 22661 53091
rect 21784 53060 22661 53088
rect 21784 53048 21790 53060
rect 22649 53057 22661 53060
rect 22695 53057 22707 53091
rect 24394 53088 24400 53100
rect 24355 53060 24400 53088
rect 22649 53051 22707 53057
rect 24394 53048 24400 53060
rect 24452 53048 24458 53100
rect 25424 53097 25452 53128
rect 26234 53116 26240 53128
rect 26292 53116 26298 53168
rect 25409 53091 25467 53097
rect 25409 53057 25421 53091
rect 25455 53057 25467 53091
rect 25409 53051 25467 53057
rect 25498 53048 25504 53100
rect 25556 53088 25562 53100
rect 25556 53060 25601 53088
rect 25556 53048 25562 53060
rect 19996 52952 20024 53048
rect 22370 53020 22376 53032
rect 22283 52992 22376 53020
rect 22370 52980 22376 52992
rect 22428 53020 22434 53032
rect 22554 53020 22560 53032
rect 22428 52992 22560 53020
rect 22428 52980 22434 52992
rect 22554 52980 22560 52992
rect 22612 52980 22618 53032
rect 24673 53023 24731 53029
rect 24673 52989 24685 53023
rect 24719 53020 24731 53023
rect 26326 53020 26332 53032
rect 24719 52992 26332 53020
rect 24719 52989 24731 52992
rect 24673 52983 24731 52989
rect 26326 52980 26332 52992
rect 26384 52980 26390 53032
rect 20993 52955 21051 52961
rect 20993 52952 21005 52955
rect 19996 52924 21005 52952
rect 20993 52921 21005 52924
rect 21039 52921 21051 52955
rect 20993 52915 21051 52921
rect 21726 52912 21732 52964
rect 21784 52952 21790 52964
rect 24026 52952 24032 52964
rect 21784 52924 24032 52952
rect 21784 52912 21790 52924
rect 24026 52912 24032 52924
rect 24084 52912 24090 52964
rect 24486 52912 24492 52964
rect 24544 52952 24550 52964
rect 26436 52952 26464 53196
rect 29748 53156 29776 53196
rect 29917 53193 29929 53227
rect 29963 53224 29975 53227
rect 31846 53224 31852 53236
rect 29963 53196 31852 53224
rect 29963 53193 29975 53196
rect 29917 53187 29975 53193
rect 31846 53184 31852 53196
rect 31904 53184 31910 53236
rect 34517 53227 34575 53233
rect 34517 53193 34529 53227
rect 34563 53224 34575 53227
rect 34790 53224 34796 53236
rect 34563 53196 34796 53224
rect 34563 53193 34575 53196
rect 34517 53187 34575 53193
rect 34790 53184 34796 53196
rect 34848 53224 34854 53236
rect 35250 53224 35256 53236
rect 34848 53196 35256 53224
rect 34848 53184 34854 53196
rect 35250 53184 35256 53196
rect 35308 53224 35314 53236
rect 35713 53227 35771 53233
rect 35713 53224 35725 53227
rect 35308 53196 35725 53224
rect 35308 53184 35314 53196
rect 35713 53193 35725 53196
rect 35759 53193 35771 53227
rect 35713 53187 35771 53193
rect 35894 53184 35900 53236
rect 35952 53224 35958 53236
rect 37090 53224 37096 53236
rect 35952 53196 37096 53224
rect 35952 53184 35958 53196
rect 37090 53184 37096 53196
rect 37148 53184 37154 53236
rect 37274 53224 37280 53236
rect 37235 53196 37280 53224
rect 37274 53184 37280 53196
rect 37332 53184 37338 53236
rect 40034 53184 40040 53236
rect 40092 53224 40098 53236
rect 40865 53227 40923 53233
rect 40865 53224 40877 53227
rect 40092 53196 40877 53224
rect 40092 53184 40098 53196
rect 40865 53193 40877 53196
rect 40911 53224 40923 53227
rect 41230 53224 41236 53236
rect 40911 53196 41236 53224
rect 40911 53193 40923 53196
rect 40865 53187 40923 53193
rect 41230 53184 41236 53196
rect 41288 53184 41294 53236
rect 41509 53227 41567 53233
rect 41509 53193 41521 53227
rect 41555 53193 41567 53227
rect 41782 53224 41788 53236
rect 41743 53196 41788 53224
rect 41509 53187 41567 53193
rect 35345 53159 35403 53165
rect 29748 53128 30880 53156
rect 27617 53091 27675 53097
rect 27617 53057 27629 53091
rect 27663 53088 27675 53091
rect 28442 53088 28448 53100
rect 27663 53060 28448 53088
rect 27663 53057 27675 53060
rect 27617 53051 27675 53057
rect 28442 53048 28448 53060
rect 28500 53048 28506 53100
rect 29086 53048 29092 53100
rect 29144 53097 29150 53100
rect 29144 53091 29172 53097
rect 29160 53057 29172 53091
rect 29144 53051 29172 53057
rect 29144 53048 29150 53051
rect 28077 53023 28135 53029
rect 28077 52989 28089 53023
rect 28123 53020 28135 53023
rect 28166 53020 28172 53032
rect 28123 52992 28172 53020
rect 28123 52989 28135 52992
rect 28077 52983 28135 52989
rect 28166 52980 28172 52992
rect 28224 52980 28230 53032
rect 28261 53023 28319 53029
rect 28261 52989 28273 53023
rect 28307 52989 28319 53023
rect 28261 52983 28319 52989
rect 24544 52924 26464 52952
rect 28276 52952 28304 52983
rect 28350 52980 28356 53032
rect 28408 53020 28414 53032
rect 28997 53023 29055 53029
rect 28997 53020 29009 53023
rect 28408 52992 29009 53020
rect 28408 52980 28414 52992
rect 28997 52989 29009 52992
rect 29043 52989 29055 53023
rect 28997 52983 29055 52989
rect 29273 53023 29331 53029
rect 29273 52989 29285 53023
rect 29319 53020 29331 53023
rect 29914 53020 29920 53032
rect 29319 52992 29920 53020
rect 29319 52989 29331 52992
rect 29273 52983 29331 52989
rect 29914 52980 29920 52992
rect 29972 53020 29978 53032
rect 30742 53020 30748 53032
rect 29972 52992 30748 53020
rect 29972 52980 29978 52992
rect 30742 52980 30748 52992
rect 30800 52980 30806 53032
rect 30852 53020 30880 53128
rect 35345 53125 35357 53159
rect 35391 53156 35403 53159
rect 35526 53156 35532 53168
rect 35391 53128 35532 53156
rect 35391 53125 35403 53128
rect 35345 53119 35403 53125
rect 35526 53116 35532 53128
rect 35584 53116 35590 53168
rect 35805 53159 35863 53165
rect 35805 53125 35817 53159
rect 35851 53156 35863 53159
rect 37918 53156 37924 53168
rect 35851 53128 37924 53156
rect 35851 53125 35863 53128
rect 35805 53119 35863 53125
rect 31113 53091 31171 53097
rect 31113 53057 31125 53091
rect 31159 53088 31171 53091
rect 32490 53088 32496 53100
rect 31159 53060 32496 53088
rect 31159 53057 31171 53060
rect 31113 53051 31171 53057
rect 32490 53048 32496 53060
rect 32548 53048 32554 53100
rect 33410 53097 33416 53100
rect 33404 53051 33416 53097
rect 33468 53088 33474 53100
rect 35621 53091 35679 53097
rect 33468 53060 33504 53088
rect 33410 53048 33416 53051
rect 33468 53048 33474 53060
rect 35621 53057 35633 53091
rect 35667 53088 35679 53091
rect 35710 53088 35716 53100
rect 35667 53060 35716 53088
rect 35667 53057 35679 53060
rect 35621 53051 35679 53057
rect 35710 53048 35716 53060
rect 35768 53048 35774 53100
rect 37458 53088 37464 53100
rect 35912 53060 37320 53088
rect 37419 53060 37464 53088
rect 30852 52992 31340 53020
rect 28721 52955 28779 52961
rect 28276 52924 28396 52952
rect 24544 52912 24550 52924
rect 1394 52844 1400 52896
rect 1452 52884 1458 52896
rect 1765 52887 1823 52893
rect 1765 52884 1777 52887
rect 1452 52856 1777 52884
rect 1452 52844 1458 52856
rect 1765 52853 1777 52856
rect 1811 52853 1823 52887
rect 1765 52847 1823 52853
rect 14921 52887 14979 52893
rect 14921 52853 14933 52887
rect 14967 52884 14979 52887
rect 15194 52884 15200 52896
rect 14967 52856 15200 52884
rect 14967 52853 14979 52856
rect 14921 52847 14979 52853
rect 15194 52844 15200 52856
rect 15252 52884 15258 52896
rect 16298 52884 16304 52896
rect 15252 52856 16304 52884
rect 15252 52844 15258 52856
rect 16298 52844 16304 52856
rect 16356 52844 16362 52896
rect 19334 52884 19340 52896
rect 19295 52856 19340 52884
rect 19334 52844 19340 52856
rect 19392 52844 19398 52896
rect 22738 52844 22744 52896
rect 22796 52884 22802 52896
rect 24578 52884 24584 52896
rect 22796 52856 24584 52884
rect 22796 52844 22802 52856
rect 24578 52844 24584 52856
rect 24636 52844 24642 52896
rect 27430 52884 27436 52896
rect 27391 52856 27436 52884
rect 27430 52844 27436 52856
rect 27488 52844 27494 52896
rect 28368 52884 28396 52924
rect 28721 52921 28733 52955
rect 28767 52952 28779 52955
rect 28810 52952 28816 52964
rect 28767 52924 28816 52952
rect 28767 52921 28779 52924
rect 28721 52915 28779 52921
rect 28810 52912 28816 52924
rect 28868 52912 28874 52964
rect 29822 52884 29828 52896
rect 28368 52856 29828 52884
rect 29822 52844 29828 52856
rect 29880 52844 29886 52896
rect 30929 52887 30987 52893
rect 30929 52853 30941 52887
rect 30975 52884 30987 52887
rect 31202 52884 31208 52896
rect 30975 52856 31208 52884
rect 30975 52853 30987 52856
rect 30929 52847 30987 52853
rect 31202 52844 31208 52856
rect 31260 52844 31266 52896
rect 31312 52884 31340 52992
rect 32766 52980 32772 53032
rect 32824 53020 32830 53032
rect 33137 53023 33195 53029
rect 33137 53020 33149 53023
rect 32824 52992 33149 53020
rect 32824 52980 32830 52992
rect 33137 52989 33149 52992
rect 33183 52989 33195 53023
rect 35912 53020 35940 53060
rect 36078 53020 36084 53032
rect 33137 52983 33195 52989
rect 35452 52992 35940 53020
rect 36039 52992 36084 53020
rect 31386 52912 31392 52964
rect 31444 52952 31450 52964
rect 32674 52952 32680 52964
rect 31444 52924 32680 52952
rect 31444 52912 31450 52924
rect 32674 52912 32680 52924
rect 32732 52912 32738 52964
rect 35452 52884 35480 52992
rect 36078 52980 36084 52992
rect 36136 52980 36142 53032
rect 37292 53020 37320 53060
rect 37458 53048 37464 53060
rect 37516 53048 37522 53100
rect 37752 53097 37780 53128
rect 37918 53116 37924 53128
rect 37976 53116 37982 53168
rect 39752 53159 39810 53165
rect 39752 53125 39764 53159
rect 39798 53156 39810 53159
rect 40770 53156 40776 53168
rect 39798 53128 40776 53156
rect 39798 53125 39810 53128
rect 39752 53119 39810 53125
rect 40770 53116 40776 53128
rect 40828 53116 40834 53168
rect 41417 53159 41475 53165
rect 41417 53125 41429 53159
rect 41463 53125 41475 53159
rect 41524 53156 41552 53187
rect 41782 53184 41788 53196
rect 41840 53184 41846 53236
rect 42794 53224 42800 53236
rect 42444 53196 42800 53224
rect 42444 53165 42472 53196
rect 42794 53184 42800 53196
rect 42852 53224 42858 53236
rect 43441 53227 43499 53233
rect 43441 53224 43453 53227
rect 42852 53196 43453 53224
rect 42852 53184 42858 53196
rect 43441 53193 43453 53196
rect 43487 53193 43499 53227
rect 45554 53224 45560 53236
rect 45515 53196 45560 53224
rect 43441 53187 43499 53193
rect 45554 53184 45560 53196
rect 45612 53184 45618 53236
rect 47946 53184 47952 53236
rect 48004 53224 48010 53236
rect 48004 53196 48084 53224
rect 48004 53184 48010 53196
rect 42429 53159 42487 53165
rect 42429 53156 42441 53159
rect 41524 53128 42441 53156
rect 41417 53119 41475 53125
rect 42429 53125 42441 53128
rect 42475 53125 42487 53159
rect 42429 53119 42487 53125
rect 37737 53091 37795 53097
rect 37737 53057 37749 53091
rect 37783 53057 37795 53091
rect 39482 53088 39488 53100
rect 39443 53060 39488 53088
rect 37737 53051 37795 53057
rect 39482 53048 39488 53060
rect 39540 53048 39546 53100
rect 41314 53091 41372 53097
rect 41314 53057 41326 53091
rect 41360 53057 41372 53091
rect 41432 53088 41460 53119
rect 42886 53116 42892 53168
rect 42944 53156 42950 53168
rect 43346 53156 43352 53168
rect 42944 53128 43352 53156
rect 42944 53116 42950 53128
rect 43346 53116 43352 53128
rect 43404 53116 43410 53168
rect 46382 53156 46388 53168
rect 45480 53128 46388 53156
rect 41432 53060 41552 53088
rect 41314 53051 41372 53057
rect 37826 53020 37832 53032
rect 37292 52992 37832 53020
rect 37826 52980 37832 52992
rect 37884 52980 37890 53032
rect 41340 53020 41368 53051
rect 41414 53020 41420 53032
rect 41340 52992 41420 53020
rect 41414 52980 41420 52992
rect 41472 52980 41478 53032
rect 41524 53020 41552 53060
rect 41598 53048 41604 53100
rect 41656 53088 41662 53100
rect 41785 53091 41843 53097
rect 41785 53088 41797 53091
rect 41656 53060 41797 53088
rect 41656 53048 41662 53060
rect 41785 53057 41797 53060
rect 41831 53057 41843 53091
rect 42610 53088 42616 53100
rect 42571 53060 42616 53088
rect 41785 53051 41843 53057
rect 42610 53048 42616 53060
rect 42668 53048 42674 53100
rect 42702 53048 42708 53100
rect 42760 53088 42766 53100
rect 44174 53088 44180 53100
rect 42760 53060 44180 53088
rect 42760 53048 42766 53060
rect 44174 53048 44180 53060
rect 44232 53048 44238 53100
rect 45480 53097 45508 53128
rect 46382 53116 46388 53128
rect 46440 53116 46446 53168
rect 46477 53159 46535 53165
rect 46477 53125 46489 53159
rect 46523 53156 46535 53159
rect 46934 53156 46940 53168
rect 46523 53128 46940 53156
rect 46523 53125 46535 53128
rect 46477 53119 46535 53125
rect 46934 53116 46940 53128
rect 46992 53116 46998 53168
rect 48056 53103 48084 53196
rect 50154 53184 50160 53236
rect 50212 53224 50218 53236
rect 50249 53227 50307 53233
rect 50249 53224 50261 53227
rect 50212 53196 50261 53224
rect 50212 53184 50218 53196
rect 50249 53193 50261 53196
rect 50295 53193 50307 53227
rect 50249 53187 50307 53193
rect 50614 53184 50620 53236
rect 50672 53224 50678 53236
rect 50893 53227 50951 53233
rect 50893 53224 50905 53227
rect 50672 53196 50905 53224
rect 50672 53184 50678 53196
rect 50893 53193 50905 53196
rect 50939 53193 50951 53227
rect 50893 53187 50951 53193
rect 45465 53091 45523 53097
rect 45465 53057 45477 53091
rect 45511 53057 45523 53091
rect 45646 53088 45652 53100
rect 45607 53060 45652 53088
rect 45465 53051 45523 53057
rect 45646 53048 45652 53060
rect 45704 53048 45710 53100
rect 46198 53048 46204 53100
rect 46256 53088 46262 53100
rect 46293 53091 46351 53097
rect 46293 53088 46305 53091
rect 46256 53060 46305 53088
rect 46256 53048 46262 53060
rect 46293 53057 46305 53060
rect 46339 53057 46351 53091
rect 46293 53051 46351 53057
rect 46569 53091 46627 53097
rect 46569 53057 46581 53091
rect 46615 53057 46627 53091
rect 47854 53088 47860 53100
rect 47815 53060 47860 53088
rect 46569 53051 46627 53057
rect 42628 53020 42656 53048
rect 41524 52992 42656 53020
rect 41616 52964 41644 52992
rect 46106 52980 46112 53032
rect 46164 53020 46170 53032
rect 46584 53020 46612 53051
rect 47854 53048 47860 53060
rect 47912 53048 47918 53100
rect 47946 53094 48004 53100
rect 47946 53060 47958 53094
rect 47992 53060 48004 53094
rect 47946 53054 48004 53060
rect 48041 53097 48099 53103
rect 48041 53063 48053 53097
rect 48087 53063 48099 53097
rect 48222 53088 48228 53100
rect 48041 53057 48099 53063
rect 48183 53060 48228 53088
rect 47581 53023 47639 53029
rect 47581 53020 47593 53023
rect 46164 52992 47593 53020
rect 46164 52980 46170 52992
rect 47581 52989 47593 52992
rect 47627 52989 47639 53023
rect 47581 52983 47639 52989
rect 35526 52912 35532 52964
rect 35584 52952 35590 52964
rect 37645 52955 37703 52961
rect 37645 52952 37657 52955
rect 35584 52924 37657 52952
rect 35584 52912 35590 52924
rect 37645 52921 37657 52924
rect 37691 52921 37703 52955
rect 37645 52915 37703 52921
rect 41598 52912 41604 52964
rect 41656 52912 41662 52964
rect 42429 52955 42487 52961
rect 42429 52952 42441 52955
rect 41708 52924 42441 52952
rect 31312 52856 35480 52884
rect 35710 52844 35716 52896
rect 35768 52884 35774 52896
rect 41708 52893 41736 52924
rect 42429 52921 42441 52924
rect 42475 52921 42487 52955
rect 47955 52952 47983 53054
rect 48222 53048 48228 53060
rect 48280 53048 48286 53100
rect 48498 53048 48504 53100
rect 48556 53088 48562 53100
rect 49878 53088 49884 53100
rect 48556 53060 49884 53088
rect 48556 53048 48562 53060
rect 49878 53048 49884 53060
rect 49936 53048 49942 53100
rect 50062 53088 50068 53100
rect 50023 53060 50068 53088
rect 50062 53048 50068 53060
rect 50120 53048 50126 53100
rect 50706 53088 50712 53100
rect 50667 53060 50712 53088
rect 50706 53048 50712 53060
rect 50764 53048 50770 53100
rect 48222 52952 48228 52964
rect 47955 52924 48228 52952
rect 42429 52915 42487 52921
rect 48222 52912 48228 52924
rect 48280 52912 48286 52964
rect 35989 52887 36047 52893
rect 35989 52884 36001 52887
rect 35768 52856 36001 52884
rect 35768 52844 35774 52856
rect 35989 52853 36001 52856
rect 36035 52853 36047 52887
rect 35989 52847 36047 52853
rect 41693 52887 41751 52893
rect 41693 52853 41705 52887
rect 41739 52853 41751 52887
rect 41693 52847 41751 52853
rect 46109 52887 46167 52893
rect 46109 52853 46121 52887
rect 46155 52884 46167 52887
rect 46290 52884 46296 52896
rect 46155 52856 46296 52884
rect 46155 52853 46167 52856
rect 46109 52847 46167 52853
rect 46290 52844 46296 52856
rect 46348 52844 46354 52896
rect 1104 52794 68816 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 65654 52794
rect 65706 52742 65718 52794
rect 65770 52742 65782 52794
rect 65834 52742 65846 52794
rect 65898 52742 65910 52794
rect 65962 52742 68816 52794
rect 1104 52720 68816 52742
rect 14090 52680 14096 52692
rect 14051 52652 14096 52680
rect 14090 52640 14096 52652
rect 14148 52640 14154 52692
rect 15286 52640 15292 52692
rect 15344 52680 15350 52692
rect 16117 52683 16175 52689
rect 16117 52680 16129 52683
rect 15344 52652 16129 52680
rect 15344 52640 15350 52652
rect 16117 52649 16129 52652
rect 16163 52649 16175 52683
rect 16117 52643 16175 52649
rect 22296 52652 23704 52680
rect 21726 52612 21732 52624
rect 21652 52584 21732 52612
rect 1394 52544 1400 52556
rect 1355 52516 1400 52544
rect 1394 52504 1400 52516
rect 1452 52504 1458 52556
rect 1854 52544 1860 52556
rect 1815 52516 1860 52544
rect 1854 52504 1860 52516
rect 1912 52504 1918 52556
rect 16574 52504 16580 52556
rect 16632 52544 16638 52556
rect 16945 52547 17003 52553
rect 16945 52544 16957 52547
rect 16632 52516 16957 52544
rect 16632 52504 16638 52516
rect 16945 52513 16957 52516
rect 16991 52513 17003 52547
rect 16945 52507 17003 52513
rect 17586 52504 17592 52556
rect 17644 52544 17650 52556
rect 18325 52547 18383 52553
rect 18325 52544 18337 52547
rect 17644 52516 18337 52544
rect 17644 52504 17650 52516
rect 18325 52513 18337 52516
rect 18371 52513 18383 52547
rect 19334 52544 19340 52556
rect 19295 52516 19340 52544
rect 18325 52507 18383 52513
rect 19334 52504 19340 52516
rect 19392 52504 19398 52556
rect 21652 52544 21680 52584
rect 21726 52572 21732 52584
rect 21784 52572 21790 52624
rect 21652 52516 21772 52544
rect 14274 52476 14280 52488
rect 14235 52448 14280 52476
rect 14274 52436 14280 52448
rect 14332 52436 14338 52488
rect 16669 52479 16727 52485
rect 16669 52445 16681 52479
rect 16715 52476 16727 52479
rect 16758 52476 16764 52488
rect 16715 52448 16764 52476
rect 16715 52445 16727 52448
rect 16669 52439 16727 52445
rect 16758 52436 16764 52448
rect 16816 52476 16822 52488
rect 17126 52476 17132 52488
rect 16816 52448 17132 52476
rect 16816 52436 16822 52448
rect 17126 52436 17132 52448
rect 17184 52436 17190 52488
rect 18046 52476 18052 52488
rect 18007 52448 18052 52476
rect 18046 52436 18052 52448
rect 18104 52436 18110 52488
rect 18138 52436 18144 52488
rect 18196 52476 18202 52488
rect 21744 52485 21772 52516
rect 21637 52479 21695 52485
rect 18196 52448 18241 52476
rect 18196 52436 18202 52448
rect 21637 52445 21649 52479
rect 21683 52445 21695 52479
rect 21637 52439 21695 52445
rect 21726 52479 21784 52485
rect 21726 52445 21738 52479
rect 21772 52445 21784 52479
rect 21726 52439 21784 52445
rect 1578 52408 1584 52420
rect 1539 52380 1584 52408
rect 1578 52368 1584 52380
rect 1636 52368 1642 52420
rect 3510 52368 3516 52420
rect 3568 52408 3574 52420
rect 3568 52380 6914 52408
rect 3568 52368 3574 52380
rect 6886 52340 6914 52380
rect 16022 52368 16028 52420
rect 16080 52408 16086 52420
rect 16080 52380 16125 52408
rect 16080 52368 16086 52380
rect 16298 52368 16304 52420
rect 16356 52408 16362 52420
rect 18322 52408 18328 52420
rect 16356 52380 18328 52408
rect 16356 52368 16362 52380
rect 18322 52368 18328 52380
rect 18380 52368 18386 52420
rect 19426 52368 19432 52420
rect 19484 52408 19490 52420
rect 19582 52411 19640 52417
rect 19582 52408 19594 52411
rect 19484 52380 19594 52408
rect 19484 52368 19490 52380
rect 19582 52377 19594 52380
rect 19628 52377 19640 52411
rect 21358 52408 21364 52420
rect 19582 52371 19640 52377
rect 19720 52380 20852 52408
rect 21319 52380 21364 52408
rect 19720 52340 19748 52380
rect 20714 52340 20720 52352
rect 6886 52312 19748 52340
rect 20675 52312 20720 52340
rect 20714 52300 20720 52312
rect 20772 52300 20778 52352
rect 20824 52340 20852 52380
rect 21358 52368 21364 52380
rect 21416 52368 21422 52420
rect 21652 52408 21680 52439
rect 21818 52436 21824 52488
rect 21876 52485 21882 52488
rect 21876 52476 21884 52485
rect 22005 52479 22063 52485
rect 21876 52448 21921 52476
rect 21876 52439 21884 52448
rect 22005 52445 22017 52479
rect 22051 52476 22063 52479
rect 22296 52476 22324 52652
rect 23676 52624 23704 52652
rect 24394 52640 24400 52692
rect 24452 52680 24458 52692
rect 28166 52680 28172 52692
rect 24452 52652 27844 52680
rect 28127 52652 28172 52680
rect 24452 52640 24458 52652
rect 23658 52572 23664 52624
rect 23716 52612 23722 52624
rect 24302 52612 24308 52624
rect 23716 52584 24308 52612
rect 23716 52572 23722 52584
rect 24302 52572 24308 52584
rect 24360 52612 24366 52624
rect 24673 52615 24731 52621
rect 24673 52612 24685 52615
rect 24360 52584 24685 52612
rect 24360 52572 24366 52584
rect 24673 52581 24685 52584
rect 24719 52581 24731 52615
rect 24673 52575 24731 52581
rect 22051 52448 22324 52476
rect 22051 52445 22063 52448
rect 22005 52439 22063 52445
rect 21876 52436 21882 52439
rect 22462 52436 22468 52488
rect 22520 52476 22526 52488
rect 23198 52476 23204 52488
rect 22520 52448 23204 52476
rect 22520 52436 22526 52448
rect 23198 52436 23204 52448
rect 23256 52436 23262 52488
rect 24210 52436 24216 52488
rect 24268 52476 24274 52488
rect 24486 52476 24492 52488
rect 24268 52448 24492 52476
rect 24268 52436 24274 52448
rect 24486 52436 24492 52448
rect 24544 52436 24550 52488
rect 25406 52476 25412 52488
rect 25367 52448 25412 52476
rect 25406 52436 25412 52448
rect 25464 52436 25470 52488
rect 26786 52476 26792 52488
rect 26747 52448 26792 52476
rect 26786 52436 26792 52448
rect 26844 52436 26850 52488
rect 27056 52479 27114 52485
rect 27056 52445 27068 52479
rect 27102 52476 27114 52479
rect 27430 52476 27436 52488
rect 27102 52448 27436 52476
rect 27102 52445 27114 52448
rect 27056 52439 27114 52445
rect 27430 52436 27436 52448
rect 27488 52436 27494 52488
rect 27816 52476 27844 52652
rect 28166 52640 28172 52652
rect 28224 52640 28230 52692
rect 28442 52640 28448 52692
rect 28500 52680 28506 52692
rect 28997 52683 29055 52689
rect 28997 52680 29009 52683
rect 28500 52652 29009 52680
rect 28500 52640 28506 52652
rect 28997 52649 29009 52652
rect 29043 52649 29055 52683
rect 28997 52643 29055 52649
rect 29086 52640 29092 52692
rect 29144 52680 29150 52692
rect 29638 52680 29644 52692
rect 29144 52652 29644 52680
rect 29144 52640 29150 52652
rect 29638 52640 29644 52652
rect 29696 52680 29702 52692
rect 29733 52683 29791 52689
rect 29733 52680 29745 52683
rect 29696 52652 29745 52680
rect 29696 52640 29702 52652
rect 29733 52649 29745 52652
rect 29779 52649 29791 52683
rect 31386 52680 31392 52692
rect 29733 52643 29791 52649
rect 29840 52652 31392 52680
rect 28184 52544 28212 52640
rect 28629 52547 28687 52553
rect 28629 52544 28641 52547
rect 28184 52516 28641 52544
rect 28629 52513 28641 52516
rect 28675 52513 28687 52547
rect 29840 52544 29868 52652
rect 31386 52640 31392 52652
rect 31444 52640 31450 52692
rect 33410 52640 33416 52692
rect 33468 52680 33474 52692
rect 33597 52683 33655 52689
rect 33597 52680 33609 52683
rect 33468 52652 33609 52680
rect 33468 52640 33474 52652
rect 33597 52649 33609 52652
rect 33643 52649 33655 52683
rect 33597 52643 33655 52649
rect 35437 52683 35495 52689
rect 35437 52649 35449 52683
rect 35483 52680 35495 52683
rect 36630 52680 36636 52692
rect 35483 52652 36636 52680
rect 35483 52649 35495 52652
rect 35437 52643 35495 52649
rect 36630 52640 36636 52652
rect 36688 52640 36694 52692
rect 43714 52680 43720 52692
rect 43675 52652 43720 52680
rect 43714 52640 43720 52652
rect 43772 52640 43778 52692
rect 46198 52640 46204 52692
rect 46256 52680 46262 52692
rect 46477 52683 46535 52689
rect 46477 52680 46489 52683
rect 46256 52652 46489 52680
rect 46256 52640 46262 52652
rect 46477 52649 46489 52652
rect 46523 52680 46535 52683
rect 48958 52680 48964 52692
rect 46523 52652 48964 52680
rect 46523 52649 46535 52652
rect 46477 52643 46535 52649
rect 48958 52640 48964 52652
rect 49016 52640 49022 52692
rect 30558 52612 30564 52624
rect 30519 52584 30564 52612
rect 30558 52572 30564 52584
rect 30616 52572 30622 52624
rect 35069 52615 35127 52621
rect 35069 52581 35081 52615
rect 35115 52612 35127 52615
rect 35526 52612 35532 52624
rect 35115 52584 35532 52612
rect 35115 52581 35127 52584
rect 35069 52575 35127 52581
rect 35526 52572 35532 52584
rect 35584 52572 35590 52624
rect 35621 52615 35679 52621
rect 35621 52581 35633 52615
rect 35667 52581 35679 52615
rect 35621 52575 35679 52581
rect 35636 52544 35664 52575
rect 37274 52572 37280 52624
rect 37332 52612 37338 52624
rect 37458 52612 37464 52624
rect 37332 52584 37464 52612
rect 37332 52572 37338 52584
rect 37458 52572 37464 52584
rect 37516 52572 37522 52624
rect 45738 52572 45744 52624
rect 45796 52612 45802 52624
rect 46661 52615 46719 52621
rect 46661 52612 46673 52615
rect 45796 52584 46673 52612
rect 45796 52572 45802 52584
rect 46661 52581 46673 52584
rect 46707 52581 46719 52615
rect 46661 52575 46719 52581
rect 28629 52507 28687 52513
rect 28736 52516 29868 52544
rect 33796 52516 35664 52544
rect 28736 52476 28764 52516
rect 27816 52448 28764 52476
rect 28813 52479 28871 52485
rect 28813 52445 28825 52479
rect 28859 52476 28871 52479
rect 28902 52476 28908 52488
rect 28859 52448 28908 52476
rect 28859 52445 28871 52448
rect 28813 52439 28871 52445
rect 28902 52436 28908 52448
rect 28960 52436 28966 52488
rect 29546 52476 29552 52488
rect 29507 52448 29552 52476
rect 29546 52436 29552 52448
rect 29604 52436 29610 52488
rect 30374 52476 30380 52488
rect 30335 52448 30380 52476
rect 30374 52436 30380 52448
rect 30432 52436 30438 52488
rect 31110 52476 31116 52488
rect 31071 52448 31116 52476
rect 31110 52436 31116 52448
rect 31168 52436 31174 52488
rect 31202 52436 31208 52488
rect 31260 52476 31266 52488
rect 33796 52485 33824 52516
rect 42610 52504 42616 52556
rect 42668 52544 42674 52556
rect 44361 52547 44419 52553
rect 44361 52544 44373 52547
rect 42668 52516 44373 52544
rect 42668 52504 42674 52516
rect 44361 52513 44373 52516
rect 44407 52544 44419 52547
rect 45554 52544 45560 52556
rect 44407 52516 45560 52544
rect 44407 52513 44419 52516
rect 44361 52507 44419 52513
rect 45554 52504 45560 52516
rect 45612 52504 45618 52556
rect 31369 52479 31427 52485
rect 31369 52476 31381 52479
rect 31260 52448 31381 52476
rect 31260 52436 31266 52448
rect 31369 52445 31381 52448
rect 31415 52445 31427 52479
rect 31369 52439 31427 52445
rect 33781 52479 33839 52485
rect 33781 52445 33793 52479
rect 33827 52445 33839 52479
rect 46106 52476 46112 52488
rect 46067 52448 46112 52476
rect 33781 52439 33839 52445
rect 46106 52436 46112 52448
rect 46164 52436 46170 52488
rect 46477 52479 46535 52485
rect 46477 52445 46489 52479
rect 46523 52476 46535 52479
rect 46566 52476 46572 52488
rect 46523 52448 46572 52476
rect 46523 52445 46535 52448
rect 46477 52439 46535 52445
rect 46566 52436 46572 52448
rect 46624 52436 46630 52488
rect 47578 52476 47584 52488
rect 47539 52448 47584 52476
rect 47578 52436 47584 52448
rect 47636 52476 47642 52488
rect 50157 52479 50215 52485
rect 50157 52476 50169 52479
rect 47636 52448 50169 52476
rect 47636 52436 47642 52448
rect 50157 52445 50169 52448
rect 50203 52476 50215 52479
rect 50706 52476 50712 52488
rect 50203 52448 50712 52476
rect 50203 52445 50215 52448
rect 50157 52439 50215 52445
rect 50706 52436 50712 52448
rect 50764 52436 50770 52488
rect 22554 52408 22560 52420
rect 21652 52380 22560 52408
rect 22554 52368 22560 52380
rect 22612 52368 22618 52420
rect 22732 52411 22790 52417
rect 22732 52377 22744 52411
rect 22778 52408 22790 52411
rect 23658 52408 23664 52420
rect 22778 52380 23664 52408
rect 22778 52377 22790 52380
rect 22732 52371 22790 52377
rect 23658 52368 23664 52380
rect 23716 52368 23722 52420
rect 34146 52408 34152 52420
rect 23768 52380 34152 52408
rect 23768 52340 23796 52380
rect 34146 52368 34152 52380
rect 34204 52368 34210 52420
rect 35434 52408 35440 52420
rect 35395 52380 35440 52408
rect 35434 52368 35440 52380
rect 35492 52368 35498 52420
rect 42334 52368 42340 52420
rect 42392 52408 42398 52420
rect 43622 52408 43628 52420
rect 42392 52380 43628 52408
rect 42392 52368 42398 52380
rect 43622 52368 43628 52380
rect 43680 52408 43686 52420
rect 45462 52408 45468 52420
rect 43680 52380 45468 52408
rect 43680 52368 43686 52380
rect 45462 52368 45468 52380
rect 45520 52368 45526 52420
rect 45554 52368 45560 52420
rect 45612 52408 45618 52420
rect 45649 52411 45707 52417
rect 45649 52408 45661 52411
rect 45612 52380 45661 52408
rect 45612 52368 45618 52380
rect 45649 52377 45661 52380
rect 45695 52408 45707 52411
rect 47854 52408 47860 52420
rect 45695 52380 47860 52408
rect 45695 52377 45707 52380
rect 45649 52371 45707 52377
rect 47854 52368 47860 52380
rect 47912 52368 47918 52420
rect 20824 52312 23796 52340
rect 23845 52343 23903 52349
rect 23845 52309 23857 52343
rect 23891 52340 23903 52343
rect 24118 52340 24124 52352
rect 23891 52312 24124 52340
rect 23891 52309 23903 52312
rect 23845 52303 23903 52309
rect 24118 52300 24124 52312
rect 24176 52300 24182 52352
rect 25130 52300 25136 52352
rect 25188 52340 25194 52352
rect 25225 52343 25283 52349
rect 25225 52340 25237 52343
rect 25188 52312 25237 52340
rect 25188 52300 25194 52312
rect 25225 52309 25237 52312
rect 25271 52309 25283 52343
rect 25225 52303 25283 52309
rect 28258 52300 28264 52352
rect 28316 52340 28322 52352
rect 28902 52340 28908 52352
rect 28316 52312 28908 52340
rect 28316 52300 28322 52312
rect 28902 52300 28908 52312
rect 28960 52300 28966 52352
rect 32122 52300 32128 52352
rect 32180 52340 32186 52352
rect 32493 52343 32551 52349
rect 32493 52340 32505 52343
rect 32180 52312 32505 52340
rect 32180 52300 32186 52312
rect 32493 52309 32505 52312
rect 32539 52309 32551 52343
rect 32493 52303 32551 52309
rect 42886 52300 42892 52352
rect 42944 52340 42950 52352
rect 44085 52343 44143 52349
rect 44085 52340 44097 52343
rect 42944 52312 44097 52340
rect 42944 52300 42950 52312
rect 44085 52309 44097 52312
rect 44131 52309 44143 52343
rect 44085 52303 44143 52309
rect 44174 52300 44180 52352
rect 44232 52340 44238 52352
rect 46934 52340 46940 52352
rect 44232 52312 46940 52340
rect 44232 52300 44238 52312
rect 46934 52300 46940 52312
rect 46992 52300 46998 52352
rect 47578 52300 47584 52352
rect 47636 52340 47642 52352
rect 47765 52343 47823 52349
rect 47765 52340 47777 52343
rect 47636 52312 47777 52340
rect 47636 52300 47642 52312
rect 47765 52309 47777 52312
rect 47811 52309 47823 52343
rect 47765 52303 47823 52309
rect 49786 52300 49792 52352
rect 49844 52340 49850 52352
rect 50341 52343 50399 52349
rect 50341 52340 50353 52343
rect 49844 52312 50353 52340
rect 49844 52300 49850 52312
rect 50341 52309 50353 52312
rect 50387 52309 50399 52343
rect 50341 52303 50399 52309
rect 1104 52250 68816 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 68816 52250
rect 1104 52176 68816 52198
rect 1578 52096 1584 52148
rect 1636 52136 1642 52148
rect 2041 52139 2099 52145
rect 2041 52136 2053 52139
rect 1636 52108 2053 52136
rect 1636 52096 1642 52108
rect 2041 52105 2053 52108
rect 2087 52105 2099 52139
rect 2041 52099 2099 52105
rect 6886 52108 55214 52136
rect 1949 52003 2007 52009
rect 1949 51969 1961 52003
rect 1995 52000 2007 52003
rect 2038 52000 2044 52012
rect 1995 51972 2044 52000
rect 1995 51969 2007 51972
rect 1949 51963 2007 51969
rect 2038 51960 2044 51972
rect 2096 52000 2102 52012
rect 6886 52000 6914 52108
rect 19705 52071 19763 52077
rect 19705 52068 19717 52071
rect 19168 52040 19717 52068
rect 2096 51972 6914 52000
rect 14636 52003 14694 52009
rect 2096 51960 2102 51972
rect 14636 51969 14648 52003
rect 14682 52000 14694 52003
rect 15010 52000 15016 52012
rect 14682 51972 15016 52000
rect 14682 51969 14694 51972
rect 14636 51963 14694 51969
rect 15010 51960 15016 51972
rect 15068 51960 15074 52012
rect 18322 51960 18328 52012
rect 18380 52000 18386 52012
rect 18380 51972 18425 52000
rect 18380 51960 18386 51972
rect 14366 51932 14372 51944
rect 14327 51904 14372 51932
rect 14366 51892 14372 51904
rect 14424 51892 14430 51944
rect 17405 51935 17463 51941
rect 17405 51901 17417 51935
rect 17451 51901 17463 51935
rect 17405 51895 17463 51901
rect 17589 51935 17647 51941
rect 17589 51901 17601 51935
rect 17635 51932 17647 51935
rect 17635 51904 18184 51932
rect 17635 51901 17647 51904
rect 17589 51895 17647 51901
rect 17420 51864 17448 51895
rect 17954 51864 17960 51876
rect 17420 51836 17960 51864
rect 17954 51824 17960 51836
rect 18012 51824 18018 51876
rect 18049 51867 18107 51873
rect 18049 51833 18061 51867
rect 18095 51833 18107 51867
rect 18049 51827 18107 51833
rect 15746 51796 15752 51808
rect 15707 51768 15752 51796
rect 15746 51756 15752 51768
rect 15804 51756 15810 51808
rect 17862 51756 17868 51808
rect 17920 51796 17926 51808
rect 18064 51796 18092 51827
rect 17920 51768 18092 51796
rect 18156 51796 18184 51904
rect 18414 51892 18420 51944
rect 18472 51941 18478 51944
rect 18472 51935 18500 51941
rect 18488 51901 18500 51935
rect 18472 51895 18500 51901
rect 18472 51892 18478 51895
rect 18598 51892 18604 51944
rect 18656 51932 18662 51944
rect 18966 51932 18972 51944
rect 18656 51904 18972 51932
rect 18656 51892 18662 51904
rect 18966 51892 18972 51904
rect 19024 51892 19030 51944
rect 19168 51796 19196 52040
rect 19705 52037 19717 52040
rect 19751 52037 19763 52071
rect 19705 52031 19763 52037
rect 19921 52071 19979 52077
rect 19921 52037 19933 52071
rect 19967 52068 19979 52071
rect 20070 52068 20076 52080
rect 19967 52040 20076 52068
rect 19967 52037 19979 52040
rect 19921 52031 19979 52037
rect 19720 52000 19748 52031
rect 20070 52028 20076 52040
rect 20128 52068 20134 52080
rect 20346 52068 20352 52080
rect 20128 52040 20352 52068
rect 20128 52028 20134 52040
rect 20346 52028 20352 52040
rect 20404 52028 20410 52080
rect 21358 52028 21364 52080
rect 21416 52068 21422 52080
rect 22066 52071 22124 52077
rect 22066 52068 22078 52071
rect 21416 52040 22078 52068
rect 21416 52028 21422 52040
rect 22066 52037 22078 52040
rect 22112 52037 22124 52071
rect 23658 52068 23664 52080
rect 22066 52031 22124 52037
rect 22572 52040 23520 52068
rect 23619 52040 23664 52068
rect 20714 52000 20720 52012
rect 19720 51972 20720 52000
rect 20714 51960 20720 51972
rect 20772 51960 20778 52012
rect 20809 52003 20867 52009
rect 20809 51969 20821 52003
rect 20855 52000 20867 52003
rect 22572 52000 22600 52040
rect 20855 51972 22600 52000
rect 23492 52000 23520 52040
rect 23658 52028 23664 52040
rect 23716 52028 23722 52080
rect 29270 52068 29276 52080
rect 23768 52040 29276 52068
rect 23768 52000 23796 52040
rect 29270 52028 29276 52040
rect 29328 52068 29334 52080
rect 29546 52068 29552 52080
rect 29328 52040 29552 52068
rect 29328 52028 29334 52040
rect 29546 52028 29552 52040
rect 29604 52028 29610 52080
rect 32122 52068 32128 52080
rect 32083 52040 32128 52068
rect 32122 52028 32128 52040
rect 32180 52028 32186 52080
rect 32355 52037 32413 52043
rect 32355 52034 32367 52037
rect 23492 51972 23796 52000
rect 23937 52003 23995 52009
rect 20855 51969 20867 51972
rect 20809 51963 20867 51969
rect 23937 51969 23949 52003
rect 23983 51969 23995 52003
rect 23937 51963 23995 51969
rect 24029 52003 24087 52009
rect 24029 51969 24041 52003
rect 24075 51969 24087 52003
rect 24029 51963 24087 51969
rect 24121 52003 24179 52009
rect 24121 51969 24133 52003
rect 24167 51969 24179 52003
rect 24302 52000 24308 52012
rect 24263 51972 24308 52000
rect 24121 51963 24179 51969
rect 19245 51935 19303 51941
rect 19245 51901 19257 51935
rect 19291 51932 19303 51935
rect 20162 51932 20168 51944
rect 19291 51904 20168 51932
rect 19291 51901 19303 51904
rect 19245 51895 19303 51901
rect 20162 51892 20168 51904
rect 20220 51892 20226 51944
rect 21821 51935 21879 51941
rect 21821 51901 21833 51935
rect 21867 51901 21879 51935
rect 23952 51932 23980 51963
rect 21821 51895 21879 51901
rect 23860 51904 23980 51932
rect 20993 51867 21051 51873
rect 20993 51864 21005 51867
rect 19260 51836 21005 51864
rect 19260 51808 19288 51836
rect 20993 51833 21005 51836
rect 21039 51833 21051 51867
rect 20993 51827 21051 51833
rect 18156 51768 19196 51796
rect 17920 51756 17926 51768
rect 19242 51756 19248 51808
rect 19300 51756 19306 51808
rect 19886 51796 19892 51808
rect 19847 51768 19892 51796
rect 19886 51756 19892 51768
rect 19944 51756 19950 51808
rect 20070 51796 20076 51808
rect 20031 51768 20076 51796
rect 20070 51756 20076 51768
rect 20128 51756 20134 51808
rect 21836 51796 21864 51895
rect 22186 51796 22192 51808
rect 21836 51768 22192 51796
rect 22186 51756 22192 51768
rect 22244 51796 22250 51808
rect 22462 51796 22468 51808
rect 22244 51768 22468 51796
rect 22244 51756 22250 51768
rect 22462 51756 22468 51768
rect 22520 51756 22526 51808
rect 22554 51756 22560 51808
rect 22612 51796 22618 51808
rect 22922 51796 22928 51808
rect 22612 51768 22928 51796
rect 22612 51756 22618 51768
rect 22922 51756 22928 51768
rect 22980 51796 22986 51808
rect 23201 51799 23259 51805
rect 23201 51796 23213 51799
rect 22980 51768 23213 51796
rect 22980 51756 22986 51768
rect 23201 51765 23213 51768
rect 23247 51765 23259 51799
rect 23860 51796 23888 51904
rect 24041 51876 24069 51963
rect 24136 51932 24164 51963
rect 24302 51960 24308 51972
rect 24360 51960 24366 52012
rect 24854 51960 24860 52012
rect 24912 52000 24918 52012
rect 25133 52003 25191 52009
rect 25133 52000 25145 52003
rect 24912 51972 25145 52000
rect 24912 51960 24918 51972
rect 25133 51969 25145 51972
rect 25179 51969 25191 52003
rect 25133 51963 25191 51969
rect 24578 51932 24584 51944
rect 24136 51904 24584 51932
rect 24578 51892 24584 51904
rect 24636 51892 24642 51944
rect 24026 51824 24032 51876
rect 24084 51824 24090 51876
rect 25148 51864 25176 51963
rect 25314 51960 25320 52012
rect 25372 52000 25378 52012
rect 25409 52003 25467 52009
rect 25409 52000 25421 52003
rect 25372 51972 25421 52000
rect 25372 51960 25378 51972
rect 25409 51969 25421 51972
rect 25455 52000 25467 52003
rect 25498 52000 25504 52012
rect 25455 51972 25504 52000
rect 25455 51969 25467 51972
rect 25409 51963 25467 51969
rect 25498 51960 25504 51972
rect 25556 51960 25562 52012
rect 28074 52000 28080 52012
rect 28035 51972 28080 52000
rect 28074 51960 28080 51972
rect 28132 51960 28138 52012
rect 28169 52003 28227 52009
rect 28169 51969 28181 52003
rect 28215 52000 28227 52003
rect 28258 52000 28264 52012
rect 28215 51972 28264 52000
rect 28215 51969 28227 51972
rect 28169 51963 28227 51969
rect 28258 51960 28264 51972
rect 28316 51960 28322 52012
rect 29641 52003 29699 52009
rect 29641 52000 29653 52003
rect 28920 51972 29653 52000
rect 28920 51944 28948 51972
rect 29641 51969 29653 51972
rect 29687 51969 29699 52003
rect 29641 51963 29699 51969
rect 29730 51960 29736 52012
rect 29788 52000 29794 52012
rect 30929 52003 30987 52009
rect 30929 52000 30941 52003
rect 29788 51972 30941 52000
rect 29788 51960 29794 51972
rect 30929 51969 30941 51972
rect 30975 52000 30987 52003
rect 32340 52003 32367 52034
rect 32401 52003 32413 52037
rect 34790 52028 34796 52080
rect 34848 52068 34854 52080
rect 35161 52071 35219 52077
rect 35161 52068 35173 52071
rect 34848 52040 35173 52068
rect 34848 52028 34854 52040
rect 35161 52037 35173 52040
rect 35207 52037 35219 52071
rect 35161 52031 35219 52037
rect 35377 52071 35435 52077
rect 35377 52037 35389 52071
rect 35423 52068 35435 52071
rect 35986 52068 35992 52080
rect 35423 52040 35992 52068
rect 35423 52037 35435 52040
rect 35377 52031 35435 52037
rect 35986 52028 35992 52040
rect 36044 52028 36050 52080
rect 41509 52071 41567 52077
rect 41509 52037 41521 52071
rect 41555 52068 41567 52071
rect 42794 52068 42800 52080
rect 41555 52040 42800 52068
rect 41555 52037 41567 52040
rect 41509 52031 41567 52037
rect 42794 52028 42800 52040
rect 42852 52028 42858 52080
rect 45833 52071 45891 52077
rect 45833 52037 45845 52071
rect 45879 52068 45891 52071
rect 47826 52071 47884 52077
rect 47826 52068 47838 52071
rect 45879 52040 47838 52068
rect 45879 52037 45891 52040
rect 45833 52031 45891 52037
rect 47826 52037 47838 52040
rect 47872 52037 47884 52071
rect 47826 52031 47884 52037
rect 32340 52000 32413 52003
rect 30975 51997 32413 52000
rect 30975 51972 32368 51997
rect 30975 51969 30987 51972
rect 30929 51963 30987 51969
rect 37550 51960 37556 52012
rect 37608 52000 37614 52012
rect 37829 52003 37887 52009
rect 37829 52000 37841 52003
rect 37608 51972 37841 52000
rect 37608 51960 37614 51972
rect 37829 51969 37841 51972
rect 37875 51969 37887 52003
rect 37829 51963 37887 51969
rect 37918 51960 37924 52012
rect 37976 52000 37982 52012
rect 38085 52003 38143 52009
rect 38085 52000 38097 52003
rect 37976 51972 38097 52000
rect 37976 51960 37982 51972
rect 38085 51969 38097 51972
rect 38131 51969 38143 52003
rect 41230 52000 41236 52012
rect 41191 51972 41236 52000
rect 38085 51963 38143 51969
rect 41230 51960 41236 51972
rect 41288 51960 41294 52012
rect 41598 52000 41604 52012
rect 41559 51972 41604 52000
rect 41598 51960 41604 51972
rect 41656 51960 41662 52012
rect 42429 52003 42487 52009
rect 42429 51969 42441 52003
rect 42475 51969 42487 52003
rect 42429 51963 42487 51969
rect 27798 51892 27804 51944
rect 27856 51932 27862 51944
rect 28902 51932 28908 51944
rect 27856 51904 28908 51932
rect 27856 51892 27862 51904
rect 28902 51892 28908 51904
rect 28960 51892 28966 51944
rect 29362 51932 29368 51944
rect 29323 51904 29368 51932
rect 29362 51892 29368 51904
rect 29420 51892 29426 51944
rect 30653 51935 30711 51941
rect 30653 51901 30665 51935
rect 30699 51901 30711 51935
rect 30653 51895 30711 51901
rect 25498 51864 25504 51876
rect 25148 51836 25504 51864
rect 25498 51824 25504 51836
rect 25556 51824 25562 51876
rect 30668 51864 30696 51895
rect 41690 51892 41696 51944
rect 41748 51941 41754 51944
rect 41748 51935 41776 51941
rect 41764 51932 41776 51935
rect 42444 51932 42472 51963
rect 43346 51960 43352 52012
rect 43404 52000 43410 52012
rect 43714 52000 43720 52012
rect 43404 51972 43720 52000
rect 43404 51960 43410 51972
rect 43714 51960 43720 51972
rect 43772 51960 43778 52012
rect 45646 51960 45652 52012
rect 45704 52000 45710 52012
rect 46109 52003 46167 52009
rect 46109 52000 46121 52003
rect 45704 51972 46121 52000
rect 45704 51960 45710 51972
rect 46109 51969 46121 51972
rect 46155 51969 46167 52003
rect 46109 51963 46167 51969
rect 46201 52003 46259 52009
rect 46201 51969 46213 52003
rect 46247 51969 46259 52003
rect 46201 51963 46259 51969
rect 43809 51935 43867 51941
rect 43809 51932 43821 51935
rect 41764 51904 42472 51932
rect 42628 51904 43821 51932
rect 41764 51901 41776 51904
rect 41748 51895 41776 51901
rect 41748 51892 41754 51895
rect 31202 51864 31208 51876
rect 27724 51836 31208 51864
rect 24118 51796 24124 51808
rect 23860 51768 24124 51796
rect 23201 51759 23259 51765
rect 24118 51756 24124 51768
rect 24176 51756 24182 51808
rect 24762 51756 24768 51808
rect 24820 51796 24826 51808
rect 27724 51796 27752 51836
rect 31202 51824 31208 51836
rect 31260 51824 31266 51876
rect 32490 51864 32496 51876
rect 32451 51836 32496 51864
rect 32490 51824 32496 51836
rect 32548 51824 32554 51876
rect 35526 51864 35532 51876
rect 35487 51836 35532 51864
rect 35526 51824 35532 51836
rect 35584 51824 35590 51876
rect 39209 51867 39267 51873
rect 39209 51833 39221 51867
rect 39255 51864 39267 51867
rect 41598 51864 41604 51876
rect 39255 51836 41604 51864
rect 39255 51833 39267 51836
rect 39209 51827 39267 51833
rect 24820 51768 27752 51796
rect 24820 51756 24826 51768
rect 27798 51756 27804 51808
rect 27856 51796 27862 51808
rect 28353 51799 28411 51805
rect 28353 51796 28365 51799
rect 27856 51768 28365 51796
rect 27856 51756 27862 51768
rect 28353 51765 28365 51768
rect 28399 51765 28411 51799
rect 28353 51759 28411 51765
rect 30006 51756 30012 51808
rect 30064 51796 30070 51808
rect 32309 51799 32367 51805
rect 32309 51796 32321 51799
rect 30064 51768 32321 51796
rect 30064 51756 30070 51768
rect 32309 51765 32321 51768
rect 32355 51765 32367 51799
rect 32309 51759 32367 51765
rect 35345 51799 35403 51805
rect 35345 51765 35357 51799
rect 35391 51796 35403 51799
rect 35618 51796 35624 51808
rect 35391 51768 35624 51796
rect 35391 51765 35403 51768
rect 35345 51759 35403 51765
rect 35618 51756 35624 51768
rect 35676 51756 35682 51808
rect 37642 51756 37648 51808
rect 37700 51796 37706 51808
rect 39224 51796 39252 51827
rect 41598 51824 41604 51836
rect 41656 51824 41662 51876
rect 41874 51824 41880 51876
rect 41932 51864 41938 51876
rect 41932 51836 41977 51864
rect 41932 51824 41938 51836
rect 37700 51768 39252 51796
rect 37700 51756 37706 51768
rect 41230 51756 41236 51808
rect 41288 51796 41294 51808
rect 42521 51799 42579 51805
rect 42521 51796 42533 51799
rect 41288 51768 42533 51796
rect 41288 51756 41294 51768
rect 42521 51765 42533 51768
rect 42567 51796 42579 51799
rect 42628 51796 42656 51904
rect 43809 51901 43821 51904
rect 43855 51932 43867 51935
rect 43990 51932 43996 51944
rect 43855 51904 43996 51932
rect 43855 51901 43867 51904
rect 43809 51895 43867 51901
rect 43990 51892 43996 51904
rect 44048 51892 44054 51944
rect 44082 51892 44088 51944
rect 44140 51892 44146 51944
rect 46216 51932 46244 51963
rect 46290 51960 46296 52012
rect 46348 52000 46354 52012
rect 46474 52000 46480 52012
rect 46348 51972 46393 52000
rect 46435 51972 46480 52000
rect 46348 51960 46354 51972
rect 46474 51960 46480 51972
rect 46532 51960 46538 52012
rect 47578 52000 47584 52012
rect 47539 51972 47584 52000
rect 47578 51960 47584 51972
rect 47636 51960 47642 52012
rect 49786 52000 49792 52012
rect 49747 51972 49792 52000
rect 49786 51960 49792 51972
rect 49844 51960 49850 52012
rect 50056 52003 50114 52009
rect 50056 51969 50068 52003
rect 50102 52000 50114 52003
rect 51074 52000 51080 52012
rect 50102 51972 51080 52000
rect 50102 51969 50114 51972
rect 50056 51963 50114 51969
rect 51074 51960 51080 51972
rect 51132 51960 51138 52012
rect 55186 52000 55214 52108
rect 67177 52003 67235 52009
rect 67177 52000 67189 52003
rect 55186 51972 67189 52000
rect 67177 51969 67189 51972
rect 67223 51969 67235 52003
rect 67177 51963 67235 51969
rect 46216 51904 46336 51932
rect 44100 51864 44128 51892
rect 46308 51876 46336 51904
rect 43916 51836 44128 51864
rect 42886 51796 42892 51808
rect 42567 51768 42656 51796
rect 42847 51768 42892 51796
rect 42567 51765 42579 51768
rect 42521 51759 42579 51765
rect 42886 51756 42892 51768
rect 42944 51756 42950 51808
rect 43916 51805 43944 51836
rect 46290 51824 46296 51876
rect 46348 51824 46354 51876
rect 48958 51864 48964 51876
rect 48919 51836 48964 51864
rect 48958 51824 48964 51836
rect 49016 51824 49022 51876
rect 43901 51799 43959 51805
rect 43901 51765 43913 51799
rect 43947 51765 43959 51799
rect 43901 51759 43959 51765
rect 44085 51799 44143 51805
rect 44085 51765 44097 51799
rect 44131 51796 44143 51799
rect 48222 51796 48228 51808
rect 44131 51768 48228 51796
rect 44131 51765 44143 51768
rect 44085 51759 44143 51765
rect 48222 51756 48228 51768
rect 48280 51756 48286 51808
rect 50522 51756 50528 51808
rect 50580 51796 50586 51808
rect 51169 51799 51227 51805
rect 51169 51796 51181 51799
rect 50580 51768 51181 51796
rect 50580 51756 50586 51768
rect 51169 51765 51181 51768
rect 51215 51765 51227 51799
rect 51169 51759 51227 51765
rect 66070 51756 66076 51808
rect 66128 51796 66134 51808
rect 67269 51799 67327 51805
rect 67269 51796 67281 51799
rect 66128 51768 67281 51796
rect 66128 51756 66134 51768
rect 67269 51765 67281 51768
rect 67315 51765 67327 51799
rect 67269 51759 67327 51765
rect 1104 51706 68816 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 65654 51706
rect 65706 51654 65718 51706
rect 65770 51654 65782 51706
rect 65834 51654 65846 51706
rect 65898 51654 65910 51706
rect 65962 51654 68816 51706
rect 1104 51632 68816 51654
rect 15010 51592 15016 51604
rect 14971 51564 15016 51592
rect 15010 51552 15016 51564
rect 15068 51552 15074 51604
rect 18046 51552 18052 51604
rect 18104 51592 18110 51604
rect 18141 51595 18199 51601
rect 18141 51592 18153 51595
rect 18104 51564 18153 51592
rect 18104 51552 18110 51564
rect 18141 51561 18153 51564
rect 18187 51561 18199 51595
rect 18141 51555 18199 51561
rect 19426 51552 19432 51604
rect 19484 51592 19490 51604
rect 19705 51595 19763 51601
rect 19705 51592 19717 51595
rect 19484 51564 19717 51592
rect 19484 51552 19490 51564
rect 19705 51561 19717 51564
rect 19751 51561 19763 51595
rect 26786 51592 26792 51604
rect 26747 51564 26792 51592
rect 19705 51555 19763 51561
rect 26786 51552 26792 51564
rect 26844 51552 26850 51604
rect 31389 51595 31447 51601
rect 31389 51561 31401 51595
rect 31435 51592 31447 51595
rect 37369 51595 37427 51601
rect 31435 51564 36584 51592
rect 31435 51561 31447 51564
rect 31389 51555 31447 51561
rect 17954 51484 17960 51536
rect 18012 51524 18018 51536
rect 19242 51524 19248 51536
rect 18012 51496 19248 51524
rect 18012 51484 18018 51496
rect 19242 51484 19248 51496
rect 19300 51484 19306 51536
rect 21818 51484 21824 51536
rect 21876 51484 21882 51536
rect 26237 51527 26295 51533
rect 26237 51493 26249 51527
rect 26283 51524 26295 51527
rect 26326 51524 26332 51536
rect 26283 51496 26332 51524
rect 26283 51493 26295 51496
rect 26237 51487 26295 51493
rect 26326 51484 26332 51496
rect 26384 51524 26390 51536
rect 26384 51496 30328 51524
rect 26384 51484 26390 51496
rect 16025 51459 16083 51465
rect 16025 51456 16037 51459
rect 15212 51428 16037 51456
rect 15212 51397 15240 51428
rect 16025 51425 16037 51428
rect 16071 51425 16083 51459
rect 16025 51419 16083 51425
rect 18138 51416 18144 51468
rect 18196 51456 18202 51468
rect 20717 51459 20775 51465
rect 20717 51456 20729 51459
rect 18196 51428 20729 51456
rect 18196 51416 18202 51428
rect 20717 51425 20729 51428
rect 20763 51425 20775 51459
rect 20717 51419 20775 51425
rect 21545 51459 21603 51465
rect 21545 51425 21557 51459
rect 21591 51456 21603 51459
rect 21836 51456 21864 51484
rect 24762 51456 24768 51468
rect 21591 51428 24768 51456
rect 21591 51425 21603 51428
rect 21545 51419 21603 51425
rect 24762 51416 24768 51428
rect 24820 51416 24826 51468
rect 28074 51416 28080 51468
rect 28132 51456 28138 51468
rect 29549 51459 29607 51465
rect 29549 51456 29561 51459
rect 28132 51428 29561 51456
rect 28132 51416 28138 51428
rect 29549 51425 29561 51428
rect 29595 51425 29607 51459
rect 29549 51419 29607 51425
rect 29638 51416 29644 51468
rect 29696 51456 29702 51468
rect 30193 51459 30251 51465
rect 30193 51456 30205 51459
rect 29696 51428 30205 51456
rect 29696 51416 29702 51428
rect 30193 51425 30205 51428
rect 30239 51425 30251 51459
rect 30300 51456 30328 51496
rect 34882 51484 34888 51536
rect 34940 51524 34946 51536
rect 35986 51524 35992 51536
rect 34940 51496 35992 51524
rect 34940 51484 34946 51496
rect 35986 51484 35992 51496
rect 36044 51484 36050 51536
rect 36446 51524 36452 51536
rect 36407 51496 36452 51524
rect 36446 51484 36452 51496
rect 36504 51484 36510 51536
rect 36556 51524 36584 51564
rect 37369 51561 37381 51595
rect 37415 51592 37427 51595
rect 37918 51592 37924 51604
rect 37415 51564 37924 51592
rect 37415 51561 37427 51564
rect 37369 51555 37427 51561
rect 37918 51552 37924 51564
rect 37976 51552 37982 51604
rect 41233 51595 41291 51601
rect 41233 51561 41245 51595
rect 41279 51592 41291 51595
rect 41690 51592 41696 51604
rect 41279 51564 41696 51592
rect 41279 51561 41291 51564
rect 41233 51555 41291 51561
rect 41690 51552 41696 51564
rect 41748 51552 41754 51604
rect 41800 51564 55214 51592
rect 36556 51496 38976 51524
rect 30586 51459 30644 51465
rect 30586 51456 30598 51459
rect 30300 51428 30598 51456
rect 30193 51419 30251 51425
rect 30586 51425 30598 51428
rect 30632 51425 30644 51459
rect 30742 51456 30748 51468
rect 30703 51428 30748 51456
rect 30586 51419 30644 51425
rect 30742 51416 30748 51428
rect 30800 51416 30806 51468
rect 34422 51416 34428 51468
rect 34480 51456 34486 51468
rect 38473 51459 38531 51465
rect 38473 51456 38485 51459
rect 34480 51428 37780 51456
rect 34480 51416 34486 51428
rect 14185 51391 14243 51397
rect 14185 51357 14197 51391
rect 14231 51388 14243 51391
rect 15197 51391 15255 51397
rect 14231 51360 14780 51388
rect 14231 51357 14243 51360
rect 14185 51351 14243 51357
rect 14752 51264 14780 51360
rect 15197 51357 15209 51391
rect 15243 51357 15255 51391
rect 15746 51388 15752 51400
rect 15659 51360 15752 51388
rect 15197 51351 15255 51357
rect 15746 51348 15752 51360
rect 15804 51348 15810 51400
rect 15841 51391 15899 51397
rect 15841 51357 15853 51391
rect 15887 51388 15899 51391
rect 16574 51388 16580 51400
rect 15887 51360 16580 51388
rect 15887 51357 15899 51360
rect 15841 51351 15899 51357
rect 16574 51348 16580 51360
rect 16632 51348 16638 51400
rect 16758 51388 16764 51400
rect 16719 51360 16764 51388
rect 16758 51348 16764 51360
rect 16816 51348 16822 51400
rect 18414 51388 18420 51400
rect 16868 51360 18420 51388
rect 15764 51320 15792 51348
rect 16868 51320 16896 51360
rect 18414 51348 18420 51360
rect 18472 51348 18478 51400
rect 19889 51391 19947 51397
rect 19889 51357 19901 51391
rect 19935 51388 19947 51391
rect 20070 51388 20076 51400
rect 19935 51360 20076 51388
rect 19935 51357 19947 51360
rect 19889 51351 19947 51357
rect 20070 51348 20076 51360
rect 20128 51348 20134 51400
rect 20346 51348 20352 51400
rect 20404 51388 20410 51400
rect 25130 51397 25136 51400
rect 21821 51391 21879 51397
rect 21821 51388 21833 51391
rect 20404 51360 21833 51388
rect 20404 51348 20410 51360
rect 21821 51357 21833 51360
rect 21867 51357 21879 51391
rect 21821 51351 21879 51357
rect 23753 51391 23811 51397
rect 23753 51357 23765 51391
rect 23799 51357 23811 51391
rect 23753 51351 23811 51357
rect 23845 51391 23903 51397
rect 23845 51357 23857 51391
rect 23891 51388 23903 51391
rect 24857 51391 24915 51397
rect 24857 51388 24869 51391
rect 23891 51360 24869 51388
rect 23891 51357 23903 51360
rect 23845 51351 23903 51357
rect 24857 51357 24869 51360
rect 24903 51357 24915 51391
rect 25124 51388 25136 51397
rect 25091 51360 25136 51388
rect 24857 51351 24915 51357
rect 25124 51351 25136 51360
rect 15764 51292 16896 51320
rect 17028 51323 17086 51329
rect 17028 51289 17040 51323
rect 17074 51320 17086 51323
rect 17402 51320 17408 51332
rect 17074 51292 17408 51320
rect 17074 51289 17086 51292
rect 17028 51283 17086 51289
rect 17402 51280 17408 51292
rect 17460 51280 17466 51332
rect 20530 51320 20536 51332
rect 20491 51292 20536 51320
rect 20530 51280 20536 51292
rect 20588 51280 20594 51332
rect 23768 51320 23796 51351
rect 25130 51348 25136 51351
rect 25188 51348 25194 51400
rect 26234 51348 26240 51400
rect 26292 51388 26298 51400
rect 26697 51391 26755 51397
rect 26697 51388 26709 51391
rect 26292 51360 26709 51388
rect 26292 51348 26298 51360
rect 26697 51357 26709 51360
rect 26743 51357 26755 51391
rect 27982 51388 27988 51400
rect 27943 51360 27988 51388
rect 26697 51351 26755 51357
rect 27982 51348 27988 51360
rect 28040 51348 28046 51400
rect 28258 51388 28264 51400
rect 28219 51360 28264 51388
rect 28258 51348 28264 51360
rect 28316 51348 28322 51400
rect 29733 51391 29791 51397
rect 29733 51357 29745 51391
rect 29779 51357 29791 51391
rect 29733 51351 29791 51357
rect 24946 51320 24952 51332
rect 23768 51292 24952 51320
rect 24946 51280 24952 51292
rect 25004 51280 25010 51332
rect 13814 51212 13820 51264
rect 13872 51252 13878 51264
rect 14369 51255 14427 51261
rect 14369 51252 14381 51255
rect 13872 51224 14381 51252
rect 13872 51212 13878 51224
rect 14369 51221 14381 51224
rect 14415 51252 14427 51255
rect 14642 51252 14648 51264
rect 14415 51224 14648 51252
rect 14415 51221 14427 51224
rect 14369 51215 14427 51221
rect 14642 51212 14648 51224
rect 14700 51212 14706 51264
rect 14734 51212 14740 51264
rect 14792 51252 14798 51264
rect 24394 51252 24400 51264
rect 14792 51224 24400 51252
rect 14792 51212 14798 51224
rect 24394 51212 24400 51224
rect 24452 51212 24458 51264
rect 29748 51252 29776 51351
rect 30466 51348 30472 51400
rect 30524 51388 30530 51400
rect 30524 51360 30569 51388
rect 30524 51348 30530 51360
rect 32030 51348 32036 51400
rect 32088 51388 32094 51400
rect 32766 51388 32772 51400
rect 32088 51360 32772 51388
rect 32088 51348 32094 51360
rect 32766 51348 32772 51360
rect 32824 51348 32830 51400
rect 34698 51388 34704 51400
rect 34659 51360 34704 51388
rect 34698 51348 34704 51360
rect 34756 51348 34762 51400
rect 34882 51388 34888 51400
rect 34843 51360 34888 51388
rect 34882 51348 34888 51360
rect 34940 51348 34946 51400
rect 35618 51348 35624 51400
rect 35676 51388 35682 51400
rect 35713 51391 35771 51397
rect 35713 51388 35725 51391
rect 35676 51360 35725 51388
rect 35676 51348 35682 51360
rect 35713 51357 35725 51360
rect 35759 51357 35771 51391
rect 35713 51351 35771 51357
rect 35802 51348 35808 51400
rect 35860 51388 35866 51400
rect 35860 51360 35905 51388
rect 35860 51348 35866 51360
rect 36354 51348 36360 51400
rect 36412 51388 36418 51400
rect 36449 51391 36507 51397
rect 36449 51388 36461 51391
rect 36412 51360 36461 51388
rect 36412 51348 36418 51360
rect 36449 51357 36461 51360
rect 36495 51357 36507 51391
rect 36722 51388 36728 51400
rect 36683 51360 36728 51388
rect 36449 51351 36507 51357
rect 36722 51348 36728 51360
rect 36780 51348 36786 51400
rect 37642 51388 37648 51400
rect 37603 51360 37648 51388
rect 37642 51348 37648 51360
rect 37700 51348 37706 51400
rect 37752 51397 37780 51428
rect 37844 51428 38485 51456
rect 37844 51397 37872 51428
rect 38473 51425 38485 51428
rect 38519 51425 38531 51459
rect 38473 51419 38531 51425
rect 37737 51391 37795 51397
rect 37737 51357 37749 51391
rect 37783 51357 37795 51391
rect 37737 51351 37795 51357
rect 37829 51391 37887 51397
rect 37829 51357 37841 51391
rect 37875 51357 37887 51391
rect 37829 51351 37887 51357
rect 38013 51391 38071 51397
rect 38013 51357 38025 51391
rect 38059 51357 38071 51391
rect 38654 51388 38660 51400
rect 38615 51360 38660 51388
rect 38013 51351 38071 51357
rect 32122 51320 32128 51332
rect 31726 51292 32128 51320
rect 31726 51252 31754 51292
rect 32122 51280 32128 51292
rect 32180 51280 32186 51332
rect 33036 51323 33094 51329
rect 33036 51289 33048 51323
rect 33082 51320 33094 51323
rect 34793 51323 34851 51329
rect 34793 51320 34805 51323
rect 33082 51292 34805 51320
rect 33082 51289 33094 51292
rect 33036 51283 33094 51289
rect 34793 51289 34805 51292
rect 34839 51289 34851 51323
rect 34793 51283 34851 51289
rect 35437 51323 35495 51329
rect 35437 51289 35449 51323
rect 35483 51320 35495 51323
rect 36078 51320 36084 51332
rect 35483 51292 36084 51320
rect 35483 51289 35495 51292
rect 35437 51283 35495 51289
rect 34146 51252 34152 51264
rect 29748 51224 31754 51252
rect 34059 51224 34152 51252
rect 34146 51212 34152 51224
rect 34204 51252 34210 51264
rect 35452 51252 35480 51283
rect 36078 51280 36084 51292
rect 36136 51280 36142 51332
rect 37090 51280 37096 51332
rect 37148 51320 37154 51332
rect 38028 51320 38056 51351
rect 38654 51348 38660 51360
rect 38712 51348 38718 51400
rect 38838 51388 38844 51400
rect 38799 51360 38844 51388
rect 38838 51348 38844 51360
rect 38896 51348 38902 51400
rect 38948 51397 38976 51496
rect 41598 51484 41604 51536
rect 41656 51524 41662 51536
rect 41800 51524 41828 51564
rect 51074 51524 51080 51536
rect 41656 51496 41828 51524
rect 42168 51496 42656 51524
rect 51035 51496 51080 51524
rect 41656 51484 41662 51496
rect 38933 51391 38991 51397
rect 38933 51357 38945 51391
rect 38979 51357 38991 51391
rect 38933 51351 38991 51357
rect 39853 51391 39911 51397
rect 39853 51357 39865 51391
rect 39899 51357 39911 51391
rect 39853 51351 39911 51357
rect 40120 51391 40178 51397
rect 40120 51357 40132 51391
rect 40166 51388 40178 51391
rect 42168 51388 42196 51496
rect 42518 51456 42524 51468
rect 42479 51428 42524 51456
rect 42518 51416 42524 51428
rect 42576 51416 42582 51468
rect 42628 51456 42656 51496
rect 51074 51484 51080 51496
rect 51132 51484 51138 51536
rect 43898 51456 43904 51468
rect 42628 51428 43904 51456
rect 43898 51416 43904 51428
rect 43956 51416 43962 51468
rect 49053 51459 49111 51465
rect 49053 51425 49065 51459
rect 49099 51456 49111 51459
rect 50062 51456 50068 51468
rect 49099 51428 50068 51456
rect 49099 51425 49111 51428
rect 49053 51419 49111 51425
rect 50062 51416 50068 51428
rect 50120 51416 50126 51468
rect 50249 51459 50307 51465
rect 50249 51425 50261 51459
rect 50295 51456 50307 51459
rect 50522 51456 50528 51468
rect 50295 51428 50528 51456
rect 50295 51425 50307 51428
rect 50249 51419 50307 51425
rect 50522 51416 50528 51428
rect 50580 51416 50586 51468
rect 55186 51456 55214 51564
rect 66257 51459 66315 51465
rect 66257 51456 66269 51459
rect 55186 51428 66269 51456
rect 66257 51425 66269 51428
rect 66303 51425 66315 51459
rect 66257 51419 66315 51425
rect 42334 51388 42340 51400
rect 40166 51360 42196 51388
rect 42295 51360 42340 51388
rect 40166 51357 40178 51360
rect 40120 51351 40178 51357
rect 39868 51320 39896 51351
rect 42334 51348 42340 51360
rect 42392 51348 42398 51400
rect 42610 51388 42616 51400
rect 42571 51360 42616 51388
rect 42610 51348 42616 51360
rect 42668 51348 42674 51400
rect 42978 51388 42984 51400
rect 42939 51360 42984 51388
rect 42978 51348 42984 51360
rect 43036 51348 43042 51400
rect 43622 51348 43628 51400
rect 43680 51388 43686 51400
rect 43717 51391 43775 51397
rect 43717 51388 43729 51391
rect 43680 51360 43729 51388
rect 43680 51348 43686 51360
rect 43717 51357 43729 51360
rect 43763 51357 43775 51391
rect 43717 51351 43775 51357
rect 43806 51348 43812 51400
rect 43864 51388 43870 51400
rect 43990 51388 43996 51400
rect 43864 51360 43909 51388
rect 43951 51360 43996 51388
rect 43864 51348 43870 51360
rect 43990 51348 43996 51360
rect 44048 51348 44054 51400
rect 44082 51348 44088 51400
rect 44140 51388 44146 51400
rect 45005 51391 45063 51397
rect 44140 51360 44185 51388
rect 44140 51348 44146 51360
rect 45005 51357 45017 51391
rect 45051 51357 45063 51391
rect 45005 51351 45063 51357
rect 37148 51292 38056 51320
rect 38764 51292 39896 51320
rect 37148 51280 37154 51292
rect 38764 51264 38792 51292
rect 41874 51280 41880 51332
rect 41932 51320 41938 51332
rect 42889 51323 42947 51329
rect 42889 51320 42901 51323
rect 41932 51292 42901 51320
rect 41932 51280 41938 51292
rect 42889 51289 42901 51292
rect 42935 51289 42947 51323
rect 42996 51320 43024 51348
rect 45020 51320 45048 51351
rect 45186 51348 45192 51400
rect 45244 51388 45250 51400
rect 45462 51388 45468 51400
rect 45244 51360 45468 51388
rect 45244 51348 45250 51360
rect 45462 51348 45468 51360
rect 45520 51348 45526 51400
rect 46017 51391 46075 51397
rect 46017 51357 46029 51391
rect 46063 51388 46075 51391
rect 46106 51388 46112 51400
rect 46063 51360 46112 51388
rect 46063 51357 46075 51360
rect 46017 51351 46075 51357
rect 46106 51348 46112 51360
rect 46164 51348 46170 51400
rect 46201 51391 46259 51397
rect 46201 51357 46213 51391
rect 46247 51388 46259 51391
rect 46566 51388 46572 51400
rect 46247 51360 46572 51388
rect 46247 51357 46259 51360
rect 46201 51351 46259 51357
rect 46566 51348 46572 51360
rect 46624 51348 46630 51400
rect 48406 51348 48412 51400
rect 48464 51388 48470 51400
rect 48777 51391 48835 51397
rect 48777 51388 48789 51391
rect 48464 51360 48789 51388
rect 48464 51348 48470 51360
rect 48777 51357 48789 51360
rect 48823 51357 48835 51391
rect 48777 51351 48835 51357
rect 50433 51391 50491 51397
rect 50433 51357 50445 51391
rect 50479 51357 50491 51391
rect 50433 51351 50491 51357
rect 50617 51391 50675 51397
rect 50617 51357 50629 51391
rect 50663 51388 50675 51391
rect 51261 51391 51319 51397
rect 51261 51388 51273 51391
rect 50663 51360 51273 51388
rect 50663 51357 50675 51360
rect 50617 51351 50675 51357
rect 51261 51357 51273 51360
rect 51307 51357 51319 51391
rect 51261 51351 51319 51357
rect 45646 51320 45652 51332
rect 42996 51292 43852 51320
rect 45020 51292 45652 51320
rect 42889 51283 42947 51289
rect 43824 51264 43852 51292
rect 45646 51280 45652 51292
rect 45704 51280 45710 51332
rect 50154 51280 50160 51332
rect 50212 51320 50218 51332
rect 50448 51320 50476 51351
rect 66438 51320 66444 51332
rect 50212 51292 50476 51320
rect 66399 51292 66444 51320
rect 50212 51280 50218 51292
rect 66438 51280 66444 51292
rect 66496 51280 66502 51332
rect 68094 51320 68100 51332
rect 68055 51292 68100 51320
rect 68094 51280 68100 51292
rect 68152 51280 68158 51332
rect 34204 51224 35480 51252
rect 34204 51212 34210 51224
rect 35526 51212 35532 51264
rect 35584 51252 35590 51264
rect 35621 51255 35679 51261
rect 35621 51252 35633 51255
rect 35584 51224 35633 51252
rect 35584 51212 35590 51224
rect 35621 51221 35633 51224
rect 35667 51252 35679 51255
rect 35710 51252 35716 51264
rect 35667 51224 35716 51252
rect 35667 51221 35679 51224
rect 35621 51215 35679 51221
rect 35710 51212 35716 51224
rect 35768 51212 35774 51264
rect 36633 51255 36691 51261
rect 36633 51221 36645 51255
rect 36679 51252 36691 51255
rect 38746 51252 38752 51264
rect 36679 51224 38752 51252
rect 36679 51221 36691 51224
rect 36633 51215 36691 51221
rect 38746 51212 38752 51224
rect 38804 51212 38810 51264
rect 43162 51212 43168 51264
rect 43220 51252 43226 51264
rect 43533 51255 43591 51261
rect 43533 51252 43545 51255
rect 43220 51224 43545 51252
rect 43220 51212 43226 51224
rect 43533 51221 43545 51224
rect 43579 51221 43591 51255
rect 43533 51215 43591 51221
rect 43806 51212 43812 51264
rect 43864 51212 43870 51264
rect 43898 51212 43904 51264
rect 43956 51252 43962 51264
rect 45097 51255 45155 51261
rect 45097 51252 45109 51255
rect 43956 51224 45109 51252
rect 43956 51212 43962 51224
rect 45097 51221 45109 51224
rect 45143 51221 45155 51255
rect 45097 51215 45155 51221
rect 45830 51212 45836 51264
rect 45888 51252 45894 51264
rect 46109 51255 46167 51261
rect 46109 51252 46121 51255
rect 45888 51224 46121 51252
rect 45888 51212 45894 51224
rect 46109 51221 46121 51224
rect 46155 51221 46167 51255
rect 46109 51215 46167 51221
rect 1104 51162 68816 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 68816 51162
rect 1104 51088 68816 51110
rect 14093 51051 14151 51057
rect 14093 51017 14105 51051
rect 14139 51048 14151 51051
rect 14366 51048 14372 51060
rect 14139 51020 14372 51048
rect 14139 51017 14151 51020
rect 14093 51011 14151 51017
rect 14366 51008 14372 51020
rect 14424 51008 14430 51060
rect 16758 51008 16764 51060
rect 16816 51048 16822 51060
rect 16853 51051 16911 51057
rect 16853 51048 16865 51051
rect 16816 51020 16865 51048
rect 16816 51008 16822 51020
rect 16853 51017 16865 51020
rect 16899 51017 16911 51051
rect 17402 51048 17408 51060
rect 17363 51020 17408 51048
rect 16853 51011 16911 51017
rect 17402 51008 17408 51020
rect 17460 51008 17466 51060
rect 20438 51008 20444 51060
rect 20496 51048 20502 51060
rect 21085 51051 21143 51057
rect 21085 51048 21097 51051
rect 20496 51020 21097 51048
rect 20496 51008 20502 51020
rect 21085 51017 21097 51020
rect 21131 51017 21143 51051
rect 21085 51011 21143 51017
rect 23661 51051 23719 51057
rect 23661 51017 23673 51051
rect 23707 51048 23719 51051
rect 23750 51048 23756 51060
rect 23707 51020 23756 51048
rect 23707 51017 23719 51020
rect 23661 51011 23719 51017
rect 23750 51008 23756 51020
rect 23808 51008 23814 51060
rect 24026 51008 24032 51060
rect 24084 51048 24090 51060
rect 24581 51051 24639 51057
rect 24581 51048 24593 51051
rect 24084 51020 24593 51048
rect 24084 51008 24090 51020
rect 24581 51017 24593 51020
rect 24627 51017 24639 51051
rect 24581 51011 24639 51017
rect 25406 51008 25412 51060
rect 25464 51048 25470 51060
rect 25685 51051 25743 51057
rect 25685 51048 25697 51051
rect 25464 51020 25697 51048
rect 25464 51008 25470 51020
rect 25685 51017 25697 51020
rect 25731 51017 25743 51051
rect 25685 51011 25743 51017
rect 28074 51008 28080 51060
rect 28132 51048 28138 51060
rect 28353 51051 28411 51057
rect 28353 51048 28365 51051
rect 28132 51020 28365 51048
rect 28132 51008 28138 51020
rect 28353 51017 28365 51020
rect 28399 51017 28411 51051
rect 28353 51011 28411 51017
rect 30466 51008 30472 51060
rect 30524 51048 30530 51060
rect 31386 51048 31392 51060
rect 30524 51020 31392 51048
rect 30524 51008 30530 51020
rect 31386 51008 31392 51020
rect 31444 51008 31450 51060
rect 31726 51020 35940 51048
rect 26326 50980 26332 50992
rect 25424 50952 26332 50980
rect 14001 50915 14059 50921
rect 14001 50881 14013 50915
rect 14047 50912 14059 50915
rect 14090 50912 14096 50924
rect 14047 50884 14096 50912
rect 14047 50881 14059 50884
rect 14001 50875 14059 50881
rect 14090 50872 14096 50884
rect 14148 50872 14154 50924
rect 14642 50912 14648 50924
rect 14603 50884 14648 50912
rect 14642 50872 14648 50884
rect 14700 50872 14706 50924
rect 16850 50912 16856 50924
rect 16763 50884 16856 50912
rect 16850 50872 16856 50884
rect 16908 50912 16914 50924
rect 17310 50912 17316 50924
rect 16908 50884 17316 50912
rect 16908 50872 16914 50884
rect 17310 50872 17316 50884
rect 17368 50872 17374 50924
rect 17586 50912 17592 50924
rect 17547 50884 17592 50912
rect 17586 50872 17592 50884
rect 17644 50872 17650 50924
rect 19705 50915 19763 50921
rect 19705 50881 19717 50915
rect 19751 50912 19763 50915
rect 20254 50912 20260 50924
rect 19751 50884 20260 50912
rect 19751 50881 19763 50884
rect 19705 50875 19763 50881
rect 20254 50872 20260 50884
rect 20312 50872 20318 50924
rect 20990 50912 20996 50924
rect 20951 50884 20996 50912
rect 20990 50872 20996 50884
rect 21048 50872 21054 50924
rect 23569 50915 23627 50921
rect 23569 50881 23581 50915
rect 23615 50912 23627 50915
rect 24394 50912 24400 50924
rect 23615 50884 24400 50912
rect 23615 50881 23627 50884
rect 23569 50875 23627 50881
rect 24394 50872 24400 50884
rect 24452 50872 24458 50924
rect 24489 50915 24547 50921
rect 24489 50881 24501 50915
rect 24535 50912 24547 50915
rect 24670 50912 24676 50924
rect 24535 50884 24676 50912
rect 24535 50881 24547 50884
rect 24489 50875 24547 50881
rect 24670 50872 24676 50884
rect 24728 50912 24734 50924
rect 25038 50912 25044 50924
rect 24728 50884 25044 50912
rect 24728 50872 24734 50884
rect 25038 50872 25044 50884
rect 25096 50872 25102 50924
rect 25424 50921 25452 50952
rect 26326 50940 26332 50952
rect 26384 50940 26390 50992
rect 30484 50980 30512 51008
rect 31110 50980 31116 50992
rect 29840 50952 30512 50980
rect 31071 50952 31116 50980
rect 25409 50915 25467 50921
rect 25409 50881 25421 50915
rect 25455 50881 25467 50915
rect 25409 50875 25467 50881
rect 25501 50915 25559 50921
rect 25501 50881 25513 50915
rect 25547 50881 25559 50915
rect 25501 50875 25559 50881
rect 25314 50804 25320 50856
rect 25372 50844 25378 50856
rect 25516 50844 25544 50875
rect 26234 50872 26240 50924
rect 26292 50912 26298 50924
rect 27240 50915 27298 50921
rect 26292 50884 26337 50912
rect 26292 50872 26298 50884
rect 27240 50881 27252 50915
rect 27286 50912 27298 50915
rect 27614 50912 27620 50924
rect 27286 50884 27620 50912
rect 27286 50881 27298 50884
rect 27240 50875 27298 50881
rect 27614 50872 27620 50884
rect 27672 50872 27678 50924
rect 29840 50921 29868 50952
rect 31110 50940 31116 50952
rect 31168 50940 31174 50992
rect 31202 50940 31208 50992
rect 31260 50980 31266 50992
rect 31726 50980 31754 51020
rect 31260 50952 31754 50980
rect 34425 50983 34483 50989
rect 31260 50940 31266 50952
rect 34425 50949 34437 50983
rect 34471 50980 34483 50983
rect 34698 50980 34704 50992
rect 34471 50952 34704 50980
rect 34471 50949 34483 50952
rect 34425 50943 34483 50949
rect 34698 50940 34704 50952
rect 34756 50940 34762 50992
rect 35434 50940 35440 50992
rect 35492 50980 35498 50992
rect 35802 50989 35808 50992
rect 35529 50983 35587 50989
rect 35529 50980 35541 50983
rect 35492 50952 35541 50980
rect 35492 50940 35498 50952
rect 35529 50949 35541 50952
rect 35575 50949 35587 50983
rect 35529 50943 35587 50949
rect 35745 50983 35808 50989
rect 35745 50949 35757 50983
rect 35791 50949 35808 50983
rect 35745 50943 35808 50949
rect 35802 50940 35808 50943
rect 35860 50940 35866 50992
rect 35912 50980 35940 51020
rect 36814 51008 36820 51060
rect 36872 51048 36878 51060
rect 46382 51048 46388 51060
rect 36872 51020 37964 51048
rect 46343 51020 46388 51048
rect 36872 51008 36878 51020
rect 35912 50952 37872 50980
rect 29825 50915 29883 50921
rect 29825 50881 29837 50915
rect 29871 50881 29883 50915
rect 29825 50875 29883 50881
rect 29917 50915 29975 50921
rect 29917 50881 29929 50915
rect 29963 50881 29975 50915
rect 29917 50875 29975 50881
rect 25372 50816 25544 50844
rect 26421 50847 26479 50853
rect 25372 50804 25378 50816
rect 26421 50813 26433 50847
rect 26467 50844 26479 50847
rect 26973 50847 27031 50853
rect 26973 50844 26985 50847
rect 26467 50816 26985 50844
rect 26467 50813 26479 50816
rect 26421 50807 26479 50813
rect 26973 50813 26985 50816
rect 27019 50813 27031 50847
rect 26973 50807 27031 50813
rect 28902 50804 28908 50856
rect 28960 50844 28966 50856
rect 29932 50844 29960 50875
rect 30558 50872 30564 50924
rect 30616 50912 30622 50924
rect 30837 50915 30895 50921
rect 30837 50912 30849 50915
rect 30616 50884 30849 50912
rect 30616 50872 30622 50884
rect 30837 50881 30849 50884
rect 30883 50881 30895 50915
rect 34146 50912 34152 50924
rect 34107 50884 34152 50912
rect 30837 50875 30895 50881
rect 34146 50872 34152 50884
rect 34204 50872 34210 50924
rect 36449 50915 36507 50921
rect 34256 50884 34560 50912
rect 34256 50844 34284 50884
rect 34422 50844 34428 50856
rect 28960 50816 29960 50844
rect 31726 50816 34284 50844
rect 34383 50816 34428 50844
rect 28960 50804 28966 50816
rect 29546 50736 29552 50788
rect 29604 50776 29610 50788
rect 29604 50748 31432 50776
rect 29604 50736 29610 50748
rect 14274 50668 14280 50720
rect 14332 50708 14338 50720
rect 14737 50711 14795 50717
rect 14737 50708 14749 50711
rect 14332 50680 14749 50708
rect 14332 50668 14338 50680
rect 14737 50677 14749 50680
rect 14783 50677 14795 50711
rect 19518 50708 19524 50720
rect 19479 50680 19524 50708
rect 14737 50671 14795 50677
rect 19518 50668 19524 50680
rect 19576 50668 19582 50720
rect 30101 50711 30159 50717
rect 30101 50677 30113 50711
rect 30147 50708 30159 50711
rect 31294 50708 31300 50720
rect 30147 50680 31300 50708
rect 30147 50677 30159 50680
rect 30101 50671 30159 50677
rect 31294 50668 31300 50680
rect 31352 50668 31358 50720
rect 31404 50708 31432 50748
rect 31726 50708 31754 50816
rect 34422 50804 34428 50816
rect 34480 50804 34486 50856
rect 34532 50844 34560 50884
rect 36449 50881 36461 50915
rect 36495 50912 36507 50915
rect 36538 50912 36544 50924
rect 36495 50884 36544 50912
rect 36495 50881 36507 50884
rect 36449 50875 36507 50881
rect 36538 50872 36544 50884
rect 36596 50912 36602 50924
rect 37737 50915 37795 50921
rect 37737 50912 37749 50915
rect 36596 50884 37749 50912
rect 36596 50872 36602 50884
rect 37737 50881 37749 50884
rect 37783 50881 37795 50915
rect 37737 50875 37795 50881
rect 37844 50844 37872 50952
rect 37936 50912 37964 51020
rect 46382 51008 46388 51020
rect 46440 51008 46446 51060
rect 46477 51051 46535 51057
rect 46477 51017 46489 51051
rect 46523 51048 46535 51051
rect 46658 51048 46664 51060
rect 46523 51020 46664 51048
rect 46523 51017 46535 51020
rect 46477 51011 46535 51017
rect 46658 51008 46664 51020
rect 46716 51008 46722 51060
rect 66438 51048 66444 51060
rect 66399 51020 66444 51048
rect 66438 51008 66444 51020
rect 66496 51008 66502 51060
rect 46109 50983 46167 50989
rect 46109 50980 46121 50983
rect 38672 50952 46121 50980
rect 38470 50912 38476 50924
rect 37936 50884 38476 50912
rect 38470 50872 38476 50884
rect 38528 50910 38534 50924
rect 38565 50915 38623 50921
rect 38565 50910 38577 50915
rect 38528 50882 38577 50910
rect 38528 50872 38534 50882
rect 38565 50881 38577 50882
rect 38611 50881 38623 50915
rect 38565 50875 38623 50881
rect 38672 50844 38700 50952
rect 46109 50949 46121 50952
rect 46155 50949 46167 50983
rect 46290 50980 46296 50992
rect 46251 50952 46296 50980
rect 46109 50943 46167 50949
rect 46290 50940 46296 50952
rect 46348 50940 46354 50992
rect 39482 50912 39488 50924
rect 39443 50884 39488 50912
rect 39482 50872 39488 50884
rect 39540 50872 39546 50924
rect 40488 50915 40546 50921
rect 40488 50881 40500 50915
rect 40534 50912 40546 50915
rect 41046 50912 41052 50924
rect 40534 50884 41052 50912
rect 40534 50881 40546 50884
rect 40488 50875 40546 50881
rect 41046 50872 41052 50884
rect 41104 50872 41110 50924
rect 43622 50872 43628 50924
rect 43680 50912 43686 50924
rect 43717 50915 43775 50921
rect 43717 50912 43729 50915
rect 43680 50884 43729 50912
rect 43680 50872 43686 50884
rect 43717 50881 43729 50884
rect 43763 50881 43775 50915
rect 43898 50912 43904 50924
rect 43859 50884 43904 50912
rect 43717 50875 43775 50881
rect 43898 50872 43904 50884
rect 43956 50912 43962 50924
rect 44082 50912 44088 50924
rect 43956 50884 44088 50912
rect 43956 50872 43962 50884
rect 44082 50872 44088 50884
rect 44140 50872 44146 50924
rect 45097 50915 45155 50921
rect 45097 50881 45109 50915
rect 45143 50912 45155 50915
rect 45646 50912 45652 50924
rect 45143 50884 45652 50912
rect 45143 50881 45155 50884
rect 45097 50875 45155 50881
rect 45646 50872 45652 50884
rect 45704 50912 45710 50924
rect 46661 50915 46719 50921
rect 46661 50912 46673 50915
rect 45704 50884 46673 50912
rect 45704 50872 45710 50884
rect 46661 50881 46673 50884
rect 46707 50881 46719 50915
rect 47670 50912 47676 50924
rect 47631 50884 47676 50912
rect 46661 50875 46719 50881
rect 47670 50872 47676 50884
rect 47728 50872 47734 50924
rect 48222 50872 48228 50924
rect 48280 50912 48286 50924
rect 48501 50915 48559 50921
rect 48501 50912 48513 50915
rect 48280 50884 48513 50912
rect 48280 50872 48286 50884
rect 48501 50881 48513 50884
rect 48547 50881 48559 50915
rect 49881 50915 49939 50921
rect 49881 50912 49893 50915
rect 48501 50875 48559 50881
rect 48608 50884 49893 50912
rect 34532 50816 36768 50844
rect 37844 50816 38700 50844
rect 39761 50847 39819 50853
rect 34238 50776 34244 50788
rect 34151 50748 34244 50776
rect 34238 50736 34244 50748
rect 34296 50776 34302 50788
rect 35897 50779 35955 50785
rect 35897 50776 35909 50779
rect 34296 50748 35909 50776
rect 34296 50736 34302 50748
rect 35897 50745 35909 50748
rect 35943 50745 35955 50779
rect 36630 50776 36636 50788
rect 36591 50748 36636 50776
rect 35897 50739 35955 50745
rect 36630 50736 36636 50748
rect 36688 50736 36694 50788
rect 31404 50680 31754 50708
rect 35710 50668 35716 50720
rect 35768 50708 35774 50720
rect 36740 50708 36768 50816
rect 39761 50813 39773 50847
rect 39807 50844 39819 50847
rect 40221 50847 40279 50853
rect 40221 50844 40233 50847
rect 39807 50816 40233 50844
rect 39807 50813 39819 50816
rect 39761 50807 39819 50813
rect 40221 50813 40233 50816
rect 40267 50813 40279 50847
rect 40221 50807 40279 50813
rect 42794 50804 42800 50856
rect 42852 50844 42858 50856
rect 43809 50847 43867 50853
rect 43809 50844 43821 50847
rect 42852 50816 43821 50844
rect 42852 50804 42858 50816
rect 43809 50813 43821 50816
rect 43855 50813 43867 50847
rect 43990 50844 43996 50856
rect 43951 50816 43996 50844
rect 43809 50807 43867 50813
rect 43990 50804 43996 50816
rect 44048 50804 44054 50856
rect 44821 50847 44879 50853
rect 44821 50813 44833 50847
rect 44867 50813 44879 50847
rect 44821 50807 44879 50813
rect 38010 50736 38016 50788
rect 38068 50776 38074 50788
rect 38657 50779 38715 50785
rect 38068 50748 38113 50776
rect 38068 50736 38074 50748
rect 38657 50745 38669 50779
rect 38703 50776 38715 50779
rect 38746 50776 38752 50788
rect 38703 50748 38752 50776
rect 38703 50745 38715 50748
rect 38657 50739 38715 50745
rect 38746 50736 38752 50748
rect 38804 50736 38810 50788
rect 41598 50776 41604 50788
rect 41559 50748 41604 50776
rect 41598 50736 41604 50748
rect 41656 50776 41662 50788
rect 42610 50776 42616 50788
rect 41656 50748 42616 50776
rect 41656 50736 41662 50748
rect 42610 50736 42616 50748
rect 42668 50736 42674 50788
rect 43533 50779 43591 50785
rect 43533 50745 43545 50779
rect 43579 50776 43591 50779
rect 44836 50776 44864 50807
rect 47026 50804 47032 50856
rect 47084 50844 47090 50856
rect 48406 50844 48412 50856
rect 47084 50816 48412 50844
rect 47084 50804 47090 50816
rect 48406 50804 48412 50816
rect 48464 50844 48470 50856
rect 48608 50844 48636 50884
rect 49881 50881 49893 50884
rect 49927 50881 49939 50915
rect 50154 50912 50160 50924
rect 50115 50884 50160 50912
rect 49881 50875 49939 50881
rect 50154 50872 50160 50884
rect 50212 50912 50218 50924
rect 51445 50915 51503 50921
rect 51445 50912 51457 50915
rect 50212 50884 51457 50912
rect 50212 50872 50218 50884
rect 51445 50881 51457 50884
rect 51491 50912 51503 50915
rect 51534 50912 51540 50924
rect 51491 50884 51540 50912
rect 51491 50881 51503 50884
rect 51445 50875 51503 50881
rect 51534 50872 51540 50884
rect 51592 50872 51598 50924
rect 51629 50915 51687 50921
rect 51629 50881 51641 50915
rect 51675 50912 51687 50915
rect 52917 50915 52975 50921
rect 52917 50912 52929 50915
rect 51675 50884 52929 50912
rect 51675 50881 51687 50884
rect 51629 50875 51687 50881
rect 52917 50881 52929 50884
rect 52963 50881 52975 50915
rect 52917 50875 52975 50881
rect 66349 50915 66407 50921
rect 66349 50881 66361 50915
rect 66395 50912 66407 50915
rect 66806 50912 66812 50924
rect 66395 50884 66812 50912
rect 66395 50881 66407 50884
rect 66349 50875 66407 50881
rect 66806 50872 66812 50884
rect 66864 50872 66870 50924
rect 48774 50844 48780 50856
rect 48464 50816 48636 50844
rect 48735 50816 48780 50844
rect 48464 50804 48470 50816
rect 48774 50804 48780 50816
rect 48832 50804 48838 50856
rect 50982 50804 50988 50856
rect 51040 50844 51046 50856
rect 51261 50847 51319 50853
rect 51261 50844 51273 50847
rect 51040 50816 51273 50844
rect 51040 50804 51046 50816
rect 51261 50813 51273 50816
rect 51307 50813 51319 50847
rect 51261 50807 51319 50813
rect 46198 50776 46204 50788
rect 43579 50748 46204 50776
rect 43579 50745 43591 50748
rect 43533 50739 43591 50745
rect 46198 50736 46204 50748
rect 46256 50776 46262 50788
rect 47118 50776 47124 50788
rect 46256 50748 47124 50776
rect 46256 50736 46262 50748
rect 47118 50736 47124 50748
rect 47176 50736 47182 50788
rect 43438 50708 43444 50720
rect 35768 50680 35813 50708
rect 36740 50680 43444 50708
rect 35768 50668 35774 50680
rect 43438 50668 43444 50680
rect 43496 50668 43502 50720
rect 47302 50668 47308 50720
rect 47360 50708 47366 50720
rect 47581 50711 47639 50717
rect 47581 50708 47593 50711
rect 47360 50680 47593 50708
rect 47360 50668 47366 50680
rect 47581 50677 47593 50680
rect 47627 50677 47639 50711
rect 48590 50708 48596 50720
rect 48551 50680 48596 50708
rect 47581 50671 47639 50677
rect 48590 50668 48596 50680
rect 48648 50668 48654 50720
rect 49050 50708 49056 50720
rect 49011 50680 49056 50708
rect 49050 50668 49056 50680
rect 49108 50668 49114 50720
rect 52730 50708 52736 50720
rect 52691 50680 52736 50708
rect 52730 50668 52736 50680
rect 52788 50668 52794 50720
rect 1104 50618 68816 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 65654 50618
rect 65706 50566 65718 50618
rect 65770 50566 65782 50618
rect 65834 50566 65846 50618
rect 65898 50566 65910 50618
rect 65962 50566 68816 50618
rect 1104 50544 68816 50566
rect 24394 50464 24400 50516
rect 24452 50504 24458 50516
rect 27614 50504 27620 50516
rect 24452 50476 26234 50504
rect 27575 50476 27620 50504
rect 24452 50464 24458 50476
rect 20990 50396 20996 50448
rect 21048 50436 21054 50448
rect 26206 50436 26234 50476
rect 27614 50464 27620 50476
rect 27672 50464 27678 50516
rect 32490 50504 32496 50516
rect 32451 50476 32496 50504
rect 32490 50464 32496 50476
rect 32548 50504 32554 50516
rect 36814 50504 36820 50516
rect 32548 50476 36820 50504
rect 32548 50464 32554 50476
rect 36814 50464 36820 50476
rect 36872 50464 36878 50516
rect 37090 50464 37096 50516
rect 37148 50504 37154 50516
rect 37148 50476 37780 50504
rect 37148 50464 37154 50476
rect 29730 50436 29736 50448
rect 21048 50408 24532 50436
rect 26206 50408 29736 50436
rect 21048 50396 21054 50408
rect 21100 50377 21128 50408
rect 21085 50371 21143 50377
rect 21085 50337 21097 50371
rect 21131 50337 21143 50371
rect 21085 50331 21143 50337
rect 21450 50328 21456 50380
rect 21508 50368 21514 50380
rect 21508 50340 22876 50368
rect 21508 50328 21514 50340
rect 12621 50303 12679 50309
rect 12621 50269 12633 50303
rect 12667 50300 12679 50303
rect 14090 50300 14096 50312
rect 12667 50272 14096 50300
rect 12667 50269 12679 50272
rect 12621 50263 12679 50269
rect 14090 50260 14096 50272
rect 14148 50260 14154 50312
rect 15102 50300 15108 50312
rect 15063 50272 15108 50300
rect 15102 50260 15108 50272
rect 15160 50260 15166 50312
rect 15194 50260 15200 50312
rect 15252 50300 15258 50312
rect 17037 50303 17095 50309
rect 15252 50272 15297 50300
rect 15252 50260 15258 50272
rect 17037 50269 17049 50303
rect 17083 50300 17095 50303
rect 18506 50300 18512 50312
rect 17083 50272 18512 50300
rect 17083 50269 17095 50272
rect 17037 50263 17095 50269
rect 18506 50260 18512 50272
rect 18564 50260 18570 50312
rect 19245 50303 19303 50309
rect 19245 50269 19257 50303
rect 19291 50300 19303 50303
rect 19334 50300 19340 50312
rect 19291 50272 19340 50300
rect 19291 50269 19303 50272
rect 19245 50263 19303 50269
rect 19334 50260 19340 50272
rect 19392 50260 19398 50312
rect 19518 50309 19524 50312
rect 19512 50300 19524 50309
rect 19479 50272 19524 50300
rect 19512 50263 19524 50272
rect 19518 50260 19524 50263
rect 19576 50260 19582 50312
rect 20070 50260 20076 50312
rect 20128 50300 20134 50312
rect 21361 50303 21419 50309
rect 21361 50300 21373 50303
rect 20128 50272 21373 50300
rect 20128 50260 20134 50272
rect 21361 50269 21373 50272
rect 21407 50269 21419 50303
rect 21361 50263 21419 50269
rect 22554 50260 22560 50312
rect 22612 50300 22618 50312
rect 22848 50309 22876 50340
rect 24118 50328 24124 50380
rect 24176 50368 24182 50380
rect 24397 50371 24455 50377
rect 24397 50368 24409 50371
rect 24176 50340 24409 50368
rect 24176 50328 24182 50340
rect 24397 50337 24409 50340
rect 24443 50337 24455 50371
rect 24504 50368 24532 50408
rect 29730 50396 29736 50408
rect 29788 50396 29794 50448
rect 37642 50436 37648 50448
rect 31726 50408 37648 50436
rect 24504 50340 27936 50368
rect 24397 50331 24455 50337
rect 22649 50303 22707 50309
rect 22649 50300 22661 50303
rect 22612 50272 22661 50300
rect 22612 50260 22618 50272
rect 22649 50269 22661 50272
rect 22695 50269 22707 50303
rect 22649 50263 22707 50269
rect 22741 50303 22799 50309
rect 22741 50269 22753 50303
rect 22787 50269 22799 50303
rect 22741 50263 22799 50269
rect 22833 50303 22891 50309
rect 22833 50269 22845 50303
rect 22879 50269 22891 50303
rect 22833 50263 22891 50269
rect 13814 50192 13820 50244
rect 13872 50232 13878 50244
rect 18598 50232 18604 50244
rect 13872 50204 18604 50232
rect 13872 50192 13878 50204
rect 18598 50192 18604 50204
rect 18656 50192 18662 50244
rect 22278 50232 22284 50244
rect 19904 50204 22284 50232
rect 12434 50124 12440 50176
rect 12492 50164 12498 50176
rect 12621 50167 12679 50173
rect 12621 50164 12633 50167
rect 12492 50136 12633 50164
rect 12492 50124 12498 50136
rect 12621 50133 12633 50136
rect 12667 50133 12679 50167
rect 15378 50164 15384 50176
rect 15339 50136 15384 50164
rect 12621 50127 12679 50133
rect 15378 50124 15384 50136
rect 15436 50124 15442 50176
rect 16574 50124 16580 50176
rect 16632 50164 16638 50176
rect 16853 50167 16911 50173
rect 16853 50164 16865 50167
rect 16632 50136 16865 50164
rect 16632 50124 16638 50136
rect 16853 50133 16865 50136
rect 16899 50133 16911 50167
rect 16853 50127 16911 50133
rect 17678 50124 17684 50176
rect 17736 50164 17742 50176
rect 19904 50164 19932 50204
rect 22278 50192 22284 50204
rect 22336 50192 22342 50244
rect 22756 50232 22784 50263
rect 23014 50260 23020 50312
rect 23072 50300 23078 50312
rect 23382 50300 23388 50312
rect 23072 50272 23388 50300
rect 23072 50260 23078 50272
rect 23382 50260 23388 50272
rect 23440 50260 23446 50312
rect 23474 50260 23480 50312
rect 23532 50300 23538 50312
rect 23569 50303 23627 50309
rect 23569 50300 23581 50303
rect 23532 50272 23581 50300
rect 23532 50260 23538 50272
rect 23569 50269 23581 50272
rect 23615 50269 23627 50303
rect 24026 50300 24032 50312
rect 23569 50263 23627 50269
rect 23676 50272 24032 50300
rect 23676 50232 23704 50272
rect 24026 50260 24032 50272
rect 24084 50260 24090 50312
rect 27798 50300 27804 50312
rect 27759 50272 27804 50300
rect 27798 50260 27804 50272
rect 27856 50260 27862 50312
rect 27908 50300 27936 50340
rect 27982 50328 27988 50380
rect 28040 50368 28046 50380
rect 31726 50368 31754 50408
rect 37642 50396 37648 50408
rect 37700 50396 37706 50448
rect 37752 50436 37780 50476
rect 38470 50464 38476 50516
rect 38528 50504 38534 50516
rect 40494 50504 40500 50516
rect 38528 50476 40500 50504
rect 38528 50464 38534 50476
rect 40494 50464 40500 50476
rect 40552 50464 40558 50516
rect 41046 50504 41052 50516
rect 41007 50476 41052 50504
rect 41046 50464 41052 50476
rect 41104 50464 41110 50516
rect 41417 50507 41475 50513
rect 41417 50473 41429 50507
rect 41463 50504 41475 50507
rect 41782 50504 41788 50516
rect 41463 50476 41788 50504
rect 41463 50473 41475 50476
rect 41417 50467 41475 50473
rect 41782 50464 41788 50476
rect 41840 50464 41846 50516
rect 47026 50504 47032 50516
rect 43364 50476 47032 50504
rect 43364 50436 43392 50476
rect 47026 50464 47032 50476
rect 47084 50464 47090 50516
rect 47302 50504 47308 50516
rect 47263 50476 47308 50504
rect 47302 50464 47308 50476
rect 47360 50464 47366 50516
rect 49050 50504 49056 50516
rect 47412 50476 49056 50504
rect 37752 50408 43392 50436
rect 43438 50396 43444 50448
rect 43496 50436 43502 50448
rect 45649 50439 45707 50445
rect 45649 50436 45661 50439
rect 43496 50408 45661 50436
rect 43496 50396 43502 50408
rect 45649 50405 45661 50408
rect 45695 50405 45707 50439
rect 47412 50436 47440 50476
rect 49050 50464 49056 50476
rect 49108 50464 49114 50516
rect 50062 50464 50068 50516
rect 50120 50504 50126 50516
rect 50341 50507 50399 50513
rect 50341 50504 50353 50507
rect 50120 50476 50353 50504
rect 50120 50464 50126 50476
rect 50341 50473 50353 50476
rect 50387 50504 50399 50507
rect 50982 50504 50988 50516
rect 50387 50476 50988 50504
rect 50387 50473 50399 50476
rect 50341 50467 50399 50473
rect 50982 50464 50988 50476
rect 51040 50504 51046 50516
rect 52917 50507 52975 50513
rect 52917 50504 52929 50507
rect 51040 50476 52929 50504
rect 51040 50464 51046 50476
rect 52917 50473 52929 50476
rect 52963 50473 52975 50507
rect 52917 50467 52975 50473
rect 48774 50436 48780 50448
rect 45649 50399 45707 50405
rect 47044 50408 47440 50436
rect 48148 50408 48780 50436
rect 41509 50371 41567 50377
rect 28040 50340 31754 50368
rect 33152 50340 38792 50368
rect 28040 50328 28046 50340
rect 29914 50300 29920 50312
rect 27908 50272 29920 50300
rect 29914 50260 29920 50272
rect 29972 50260 29978 50312
rect 30006 50260 30012 50312
rect 30064 50300 30070 50312
rect 30193 50303 30251 50309
rect 30193 50300 30205 50303
rect 30064 50272 30205 50300
rect 30064 50260 30070 50272
rect 30193 50269 30205 50272
rect 30239 50269 30251 50303
rect 30193 50263 30251 50269
rect 30282 50260 30288 50312
rect 30340 50300 30346 50312
rect 32309 50303 32367 50309
rect 32309 50300 32321 50303
rect 30340 50272 32321 50300
rect 30340 50260 30346 50272
rect 32309 50269 32321 50272
rect 32355 50300 32367 50303
rect 32582 50300 32588 50312
rect 32355 50272 32588 50300
rect 32355 50269 32367 50272
rect 32309 50263 32367 50269
rect 32582 50260 32588 50272
rect 32640 50260 32646 50312
rect 22756 50204 23704 50232
rect 23845 50235 23903 50241
rect 23845 50201 23857 50235
rect 23891 50232 23903 50235
rect 24581 50235 24639 50241
rect 24581 50232 24593 50235
rect 23891 50204 24593 50232
rect 23891 50201 23903 50204
rect 23845 50195 23903 50201
rect 24581 50201 24593 50204
rect 24627 50201 24639 50235
rect 24581 50195 24639 50201
rect 17736 50136 19932 50164
rect 17736 50124 17742 50136
rect 19978 50124 19984 50176
rect 20036 50164 20042 50176
rect 20625 50167 20683 50173
rect 20625 50164 20637 50167
rect 20036 50136 20637 50164
rect 20036 50124 20042 50136
rect 20625 50133 20637 50136
rect 20671 50133 20683 50167
rect 22370 50164 22376 50176
rect 22331 50136 22376 50164
rect 20625 50127 20683 50133
rect 22370 50124 22376 50136
rect 22428 50124 22434 50176
rect 24596 50164 24624 50195
rect 25866 50192 25872 50244
rect 25924 50232 25930 50244
rect 26237 50235 26295 50241
rect 26237 50232 26249 50235
rect 25924 50204 26249 50232
rect 25924 50192 25930 50204
rect 26237 50201 26249 50204
rect 26283 50201 26295 50235
rect 33152 50232 33180 50340
rect 33229 50303 33287 50309
rect 33229 50269 33241 50303
rect 33275 50300 33287 50303
rect 35161 50303 35219 50309
rect 35161 50300 35173 50303
rect 33275 50272 35173 50300
rect 33275 50269 33287 50272
rect 33229 50263 33287 50269
rect 35161 50269 35173 50272
rect 35207 50300 35219 50303
rect 36078 50300 36084 50312
rect 35207 50272 36084 50300
rect 35207 50269 35219 50272
rect 35161 50263 35219 50269
rect 36078 50260 36084 50272
rect 36136 50260 36142 50312
rect 36357 50303 36415 50309
rect 36357 50269 36369 50303
rect 36403 50300 36415 50303
rect 36538 50300 36544 50312
rect 36403 50272 36544 50300
rect 36403 50269 36415 50272
rect 36357 50263 36415 50269
rect 36538 50260 36544 50272
rect 36596 50260 36602 50312
rect 38289 50303 38347 50309
rect 38289 50269 38301 50303
rect 38335 50300 38347 50303
rect 38562 50300 38568 50312
rect 38335 50272 38568 50300
rect 38335 50269 38347 50272
rect 38289 50263 38347 50269
rect 38562 50260 38568 50272
rect 38620 50260 38626 50312
rect 38764 50309 38792 50340
rect 41509 50337 41521 50371
rect 41555 50368 41567 50371
rect 41598 50368 41604 50380
rect 41555 50340 41604 50368
rect 41555 50337 41567 50340
rect 41509 50331 41567 50337
rect 41598 50328 41604 50340
rect 41656 50328 41662 50380
rect 38749 50303 38807 50309
rect 38749 50269 38761 50303
rect 38795 50269 38807 50303
rect 38749 50263 38807 50269
rect 39666 50260 39672 50312
rect 39724 50300 39730 50312
rect 39945 50303 40003 50309
rect 39945 50300 39957 50303
rect 39724 50272 39957 50300
rect 39724 50260 39730 50272
rect 39945 50269 39957 50272
rect 39991 50269 40003 50303
rect 39945 50263 40003 50269
rect 41233 50303 41291 50309
rect 41233 50269 41245 50303
rect 41279 50300 41291 50303
rect 41322 50300 41328 50312
rect 41279 50272 41328 50300
rect 41279 50269 41291 50272
rect 41233 50263 41291 50269
rect 41322 50260 41328 50272
rect 41380 50260 41386 50312
rect 41874 50260 41880 50312
rect 41932 50300 41938 50312
rect 42426 50300 42432 50312
rect 41932 50272 42432 50300
rect 41932 50260 41938 50272
rect 42426 50260 42432 50272
rect 42484 50260 42490 50312
rect 45830 50300 45836 50312
rect 45791 50272 45836 50300
rect 45830 50260 45836 50272
rect 45888 50260 45894 50312
rect 46290 50260 46296 50312
rect 46348 50300 46354 50312
rect 47044 50309 47072 50408
rect 47118 50328 47124 50380
rect 47176 50368 47182 50380
rect 47176 50340 47221 50368
rect 47176 50328 47182 50340
rect 47029 50303 47087 50309
rect 47029 50300 47041 50303
rect 46348 50272 47041 50300
rect 46348 50260 46354 50272
rect 47029 50269 47041 50272
rect 47075 50269 47087 50303
rect 47029 50263 47087 50269
rect 47305 50303 47363 50309
rect 47305 50269 47317 50303
rect 47351 50269 47363 50303
rect 47305 50263 47363 50269
rect 26237 50195 26295 50201
rect 29840 50204 33180 50232
rect 29840 50164 29868 50204
rect 34422 50192 34428 50244
rect 34480 50232 34486 50244
rect 36630 50232 36636 50244
rect 34480 50204 36636 50232
rect 34480 50192 34486 50204
rect 36630 50192 36636 50204
rect 36688 50192 36694 50244
rect 37550 50232 37556 50244
rect 37511 50204 37556 50232
rect 37550 50192 37556 50204
rect 37608 50232 37614 50244
rect 38657 50235 38715 50241
rect 38657 50232 38669 50235
rect 37608 50204 38669 50232
rect 37608 50192 37614 50204
rect 38657 50201 38669 50204
rect 38703 50201 38715 50235
rect 44082 50232 44088 50244
rect 38657 50195 38715 50201
rect 38764 50204 44088 50232
rect 24596 50136 29868 50164
rect 29914 50124 29920 50176
rect 29972 50164 29978 50176
rect 33318 50164 33324 50176
rect 29972 50136 33324 50164
rect 29972 50124 29978 50136
rect 33318 50124 33324 50136
rect 33376 50164 33382 50176
rect 33413 50167 33471 50173
rect 33413 50164 33425 50167
rect 33376 50136 33425 50164
rect 33376 50124 33382 50136
rect 33413 50133 33425 50136
rect 33459 50133 33471 50167
rect 33413 50127 33471 50133
rect 35437 50167 35495 50173
rect 35437 50133 35449 50167
rect 35483 50164 35495 50167
rect 35710 50164 35716 50176
rect 35483 50136 35716 50164
rect 35483 50133 35495 50136
rect 35437 50127 35495 50133
rect 35710 50124 35716 50136
rect 35768 50164 35774 50176
rect 37090 50164 37096 50176
rect 35768 50136 37096 50164
rect 35768 50124 35774 50136
rect 37090 50124 37096 50136
rect 37148 50124 37154 50176
rect 37458 50124 37464 50176
rect 37516 50164 37522 50176
rect 37645 50167 37703 50173
rect 37645 50164 37657 50167
rect 37516 50136 37657 50164
rect 37516 50124 37522 50136
rect 37645 50133 37657 50136
rect 37691 50164 37703 50167
rect 37734 50164 37740 50176
rect 37691 50136 37740 50164
rect 37691 50133 37703 50136
rect 37645 50127 37703 50133
rect 37734 50124 37740 50136
rect 37792 50124 37798 50176
rect 38010 50124 38016 50176
rect 38068 50164 38074 50176
rect 38764 50164 38792 50204
rect 44082 50192 44088 50204
rect 44140 50192 44146 50244
rect 45646 50192 45652 50244
rect 45704 50232 45710 50244
rect 46201 50235 46259 50241
rect 46201 50232 46213 50235
rect 45704 50204 46213 50232
rect 45704 50192 45710 50204
rect 46201 50201 46213 50204
rect 46247 50201 46259 50235
rect 47320 50232 47348 50263
rect 47762 50260 47768 50312
rect 47820 50300 47826 50312
rect 48148 50309 48176 50408
rect 48774 50396 48780 50408
rect 48832 50436 48838 50448
rect 50709 50439 50767 50445
rect 50709 50436 50721 50439
rect 48832 50408 50721 50436
rect 48832 50396 48838 50408
rect 50709 50405 50721 50408
rect 50755 50405 50767 50439
rect 50709 50399 50767 50405
rect 48222 50328 48228 50380
rect 48280 50368 48286 50380
rect 48280 50340 48912 50368
rect 48280 50328 48286 50340
rect 48133 50303 48191 50309
rect 48133 50300 48145 50303
rect 47820 50272 48145 50300
rect 47820 50260 47826 50272
rect 48133 50269 48145 50272
rect 48179 50269 48191 50303
rect 48133 50263 48191 50269
rect 48501 50303 48559 50309
rect 48501 50269 48513 50303
rect 48547 50300 48559 50303
rect 48590 50300 48596 50312
rect 48547 50272 48596 50300
rect 48547 50269 48559 50272
rect 48501 50263 48559 50269
rect 48314 50232 48320 50244
rect 47320 50204 48320 50232
rect 46201 50195 46259 50201
rect 48314 50192 48320 50204
rect 48372 50192 48378 50244
rect 48516 50232 48544 50263
rect 48590 50260 48596 50272
rect 48648 50260 48654 50312
rect 48884 50309 48912 50340
rect 48869 50303 48927 50309
rect 48869 50269 48881 50303
rect 48915 50269 48927 50303
rect 48869 50263 48927 50269
rect 50154 50260 50160 50312
rect 50212 50300 50218 50312
rect 50341 50303 50399 50309
rect 50341 50300 50353 50303
rect 50212 50272 50353 50300
rect 50212 50260 50218 50272
rect 50341 50269 50353 50272
rect 50387 50269 50399 50303
rect 50341 50263 50399 50269
rect 50525 50303 50583 50309
rect 50525 50269 50537 50303
rect 50571 50300 50583 50303
rect 50614 50300 50620 50312
rect 50571 50272 50620 50300
rect 50571 50269 50583 50272
rect 50525 50263 50583 50269
rect 50614 50260 50620 50272
rect 50672 50260 50678 50312
rect 51350 50260 51356 50312
rect 51408 50300 51414 50312
rect 51537 50303 51595 50309
rect 51537 50300 51549 50303
rect 51408 50272 51549 50300
rect 51408 50260 51414 50272
rect 51537 50269 51549 50272
rect 51583 50269 51595 50303
rect 51537 50263 51595 50269
rect 51804 50303 51862 50309
rect 51804 50269 51816 50303
rect 51850 50300 51862 50303
rect 52730 50300 52736 50312
rect 51850 50272 52736 50300
rect 51850 50269 51862 50272
rect 51804 50263 51862 50269
rect 52730 50260 52736 50272
rect 52788 50260 52794 50312
rect 49786 50232 49792 50244
rect 48516 50204 49792 50232
rect 49786 50192 49792 50204
rect 49844 50192 49850 50244
rect 38068 50136 38792 50164
rect 40129 50167 40187 50173
rect 38068 50124 38074 50136
rect 40129 50133 40141 50167
rect 40175 50164 40187 50167
rect 41966 50164 41972 50176
rect 40175 50136 41972 50164
rect 40175 50133 40187 50136
rect 40129 50127 40187 50133
rect 41966 50124 41972 50136
rect 42024 50164 42030 50176
rect 43070 50164 43076 50176
rect 42024 50136 43076 50164
rect 42024 50124 42030 50136
rect 43070 50124 43076 50136
rect 43128 50124 43134 50176
rect 45922 50164 45928 50176
rect 45883 50136 45928 50164
rect 45922 50124 45928 50136
rect 45980 50124 45986 50176
rect 46017 50167 46075 50173
rect 46017 50133 46029 50167
rect 46063 50164 46075 50167
rect 46106 50164 46112 50176
rect 46063 50136 46112 50164
rect 46063 50133 46075 50136
rect 46017 50127 46075 50133
rect 46106 50124 46112 50136
rect 46164 50124 46170 50176
rect 47486 50164 47492 50176
rect 47447 50136 47492 50164
rect 47486 50124 47492 50136
rect 47544 50124 47550 50176
rect 48130 50164 48136 50176
rect 48091 50136 48136 50164
rect 48130 50124 48136 50136
rect 48188 50124 48194 50176
rect 1104 50074 68816 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 68816 50074
rect 1104 50000 68816 50022
rect 3510 49920 3516 49972
rect 3568 49960 3574 49972
rect 17678 49960 17684 49972
rect 3568 49932 17684 49960
rect 3568 49920 3574 49932
rect 17678 49920 17684 49932
rect 17736 49920 17742 49972
rect 19978 49960 19984 49972
rect 17788 49932 19984 49960
rect 12434 49824 12440 49836
rect 12395 49796 12440 49824
rect 12434 49784 12440 49796
rect 12492 49784 12498 49836
rect 12704 49827 12762 49833
rect 12704 49793 12716 49827
rect 12750 49824 12762 49827
rect 12986 49824 12992 49836
rect 12750 49796 12992 49824
rect 12750 49793 12762 49796
rect 12704 49787 12762 49793
rect 12986 49784 12992 49796
rect 13044 49784 13050 49836
rect 14274 49824 14280 49836
rect 14235 49796 14280 49824
rect 14274 49784 14280 49796
rect 14332 49784 14338 49836
rect 14366 49784 14372 49836
rect 14424 49824 14430 49836
rect 14533 49827 14591 49833
rect 14533 49824 14545 49827
rect 14424 49796 14545 49824
rect 14424 49784 14430 49796
rect 14533 49793 14545 49796
rect 14579 49793 14591 49827
rect 14533 49787 14591 49793
rect 15102 49784 15108 49836
rect 15160 49824 15166 49836
rect 16850 49824 16856 49836
rect 15160 49796 15608 49824
rect 16811 49796 16856 49824
rect 15160 49784 15166 49796
rect 15580 49756 15608 49796
rect 16850 49784 16856 49796
rect 16908 49784 16914 49836
rect 15580 49728 17540 49756
rect 13814 49688 13820 49700
rect 13775 49660 13820 49688
rect 13814 49648 13820 49660
rect 13872 49648 13878 49700
rect 15672 49697 15700 49728
rect 15657 49691 15715 49697
rect 15657 49657 15669 49691
rect 15703 49657 15715 49691
rect 17512 49688 17540 49728
rect 17586 49716 17592 49768
rect 17644 49756 17650 49768
rect 17788 49765 17816 49932
rect 19904 49901 19932 49932
rect 19978 49920 19984 49932
rect 20036 49920 20042 49972
rect 20254 49960 20260 49972
rect 20215 49932 20260 49960
rect 20254 49920 20260 49932
rect 20312 49920 20318 49972
rect 24946 49960 24952 49972
rect 24907 49932 24952 49960
rect 24946 49920 24952 49932
rect 25004 49920 25010 49972
rect 25130 49920 25136 49972
rect 25188 49960 25194 49972
rect 25498 49960 25504 49972
rect 25188 49932 25504 49960
rect 25188 49920 25194 49932
rect 25498 49920 25504 49932
rect 25556 49960 25562 49972
rect 25556 49932 29332 49960
rect 25556 49920 25562 49932
rect 19889 49895 19947 49901
rect 19889 49861 19901 49895
rect 19935 49861 19947 49895
rect 19889 49855 19947 49861
rect 20089 49895 20147 49901
rect 20089 49861 20101 49895
rect 20135 49892 20147 49895
rect 20135 49864 20208 49892
rect 20135 49861 20147 49864
rect 20089 49855 20147 49861
rect 18598 49784 18604 49836
rect 18656 49833 18662 49836
rect 18656 49827 18684 49833
rect 18672 49793 18684 49827
rect 20180 49824 20208 49864
rect 22278 49852 22284 49904
rect 22336 49892 22342 49904
rect 22336 49864 23888 49892
rect 22336 49852 22342 49864
rect 20254 49824 20260 49836
rect 20180 49796 20260 49824
rect 18656 49787 18684 49793
rect 18656 49784 18662 49787
rect 20254 49784 20260 49796
rect 20312 49784 20318 49836
rect 17773 49759 17831 49765
rect 17644 49728 17689 49756
rect 17644 49716 17650 49728
rect 17773 49725 17785 49759
rect 17819 49725 17831 49759
rect 18509 49759 18567 49765
rect 18509 49756 18521 49759
rect 17773 49719 17831 49725
rect 17880 49728 18521 49756
rect 17880 49688 17908 49728
rect 18509 49725 18521 49728
rect 18555 49725 18567 49759
rect 18509 49719 18567 49725
rect 18785 49759 18843 49765
rect 18785 49725 18797 49759
rect 18831 49756 18843 49759
rect 18966 49756 18972 49768
rect 18831 49728 18972 49756
rect 18831 49725 18843 49728
rect 18785 49719 18843 49725
rect 18966 49716 18972 49728
rect 19024 49716 19030 49768
rect 19429 49759 19487 49765
rect 19429 49725 19441 49759
rect 19475 49756 19487 49759
rect 20622 49756 20628 49768
rect 19475 49728 20628 49756
rect 19475 49725 19487 49728
rect 19429 49719 19487 49725
rect 20622 49716 20628 49728
rect 20680 49716 20686 49768
rect 22465 49759 22523 49765
rect 22465 49725 22477 49759
rect 22511 49725 22523 49759
rect 22465 49719 22523 49725
rect 22649 49759 22707 49765
rect 22649 49725 22661 49759
rect 22695 49756 22707 49759
rect 22830 49756 22836 49768
rect 22695 49728 22836 49756
rect 22695 49725 22707 49728
rect 22649 49719 22707 49725
rect 18230 49688 18236 49700
rect 17512 49660 17908 49688
rect 18191 49660 18236 49688
rect 15657 49651 15715 49657
rect 18230 49648 18236 49660
rect 18288 49648 18294 49700
rect 22480 49688 22508 49719
rect 22830 49716 22836 49728
rect 22888 49716 22894 49768
rect 23860 49765 23888 49864
rect 24394 49784 24400 49836
rect 24452 49824 24458 49836
rect 24765 49827 24823 49833
rect 24765 49824 24777 49827
rect 24452 49796 24777 49824
rect 24452 49784 24458 49796
rect 24765 49793 24777 49796
rect 24811 49793 24823 49827
rect 24765 49787 24823 49793
rect 26237 49827 26295 49833
rect 26237 49793 26249 49827
rect 26283 49824 26295 49827
rect 27338 49824 27344 49836
rect 26283 49796 27344 49824
rect 26283 49793 26295 49796
rect 26237 49787 26295 49793
rect 27338 49784 27344 49796
rect 27396 49784 27402 49836
rect 28813 49827 28871 49833
rect 28813 49793 28825 49827
rect 28859 49824 28871 49827
rect 29178 49824 29184 49836
rect 28859 49796 29184 49824
rect 28859 49793 28871 49796
rect 28813 49787 28871 49793
rect 29178 49784 29184 49796
rect 29236 49784 29242 49836
rect 23845 49759 23903 49765
rect 23845 49725 23857 49759
rect 23891 49725 23903 49759
rect 23845 49719 23903 49725
rect 22554 49688 22560 49700
rect 22467 49660 22560 49688
rect 22554 49648 22560 49660
rect 22612 49688 22618 49700
rect 23014 49688 23020 49700
rect 22612 49660 23020 49688
rect 22612 49648 22618 49660
rect 23014 49648 23020 49660
rect 23072 49648 23078 49700
rect 16850 49620 16856 49632
rect 16811 49592 16856 49620
rect 16850 49580 16856 49592
rect 16908 49580 16914 49632
rect 20070 49620 20076 49632
rect 20031 49592 20076 49620
rect 20070 49580 20076 49592
rect 20128 49580 20134 49632
rect 26050 49620 26056 49632
rect 26011 49592 26056 49620
rect 26050 49580 26056 49592
rect 26108 49580 26114 49632
rect 28626 49620 28632 49632
rect 28587 49592 28632 49620
rect 28626 49580 28632 49592
rect 28684 49580 28690 49632
rect 29304 49620 29332 49932
rect 32582 49920 32588 49972
rect 32640 49960 32646 49972
rect 33505 49963 33563 49969
rect 33505 49960 33517 49963
rect 32640 49932 33517 49960
rect 32640 49920 32646 49932
rect 33505 49929 33517 49932
rect 33551 49929 33563 49963
rect 36633 49963 36691 49969
rect 36633 49960 36645 49963
rect 33505 49923 33563 49929
rect 33612 49932 36645 49960
rect 33612 49892 33640 49932
rect 36633 49929 36645 49932
rect 36679 49929 36691 49963
rect 36633 49923 36691 49929
rect 37366 49920 37372 49972
rect 37424 49960 37430 49972
rect 37461 49963 37519 49969
rect 37461 49960 37473 49963
rect 37424 49932 37473 49960
rect 37424 49920 37430 49932
rect 37461 49929 37473 49932
rect 37507 49929 37519 49963
rect 37461 49923 37519 49929
rect 37642 49920 37648 49972
rect 37700 49960 37706 49972
rect 43717 49963 43775 49969
rect 43717 49960 43729 49963
rect 37700 49932 41828 49960
rect 37700 49920 37706 49932
rect 30208 49864 33640 49892
rect 34609 49895 34667 49901
rect 29365 49827 29423 49833
rect 29365 49793 29377 49827
rect 29411 49824 29423 49827
rect 30098 49824 30104 49836
rect 29411 49796 30104 49824
rect 29411 49793 29423 49796
rect 29365 49787 29423 49793
rect 30098 49784 30104 49796
rect 30156 49784 30162 49836
rect 30208 49833 30236 49864
rect 34609 49861 34621 49895
rect 34655 49892 34667 49895
rect 35253 49895 35311 49901
rect 35253 49892 35265 49895
rect 34655 49864 35265 49892
rect 34655 49861 34667 49864
rect 34609 49855 34667 49861
rect 35253 49861 35265 49864
rect 35299 49861 35311 49895
rect 35253 49855 35311 49861
rect 36078 49852 36084 49904
rect 36136 49892 36142 49904
rect 36136 49864 37504 49892
rect 36136 49852 36142 49864
rect 30193 49827 30251 49833
rect 30193 49793 30205 49827
rect 30239 49793 30251 49827
rect 30193 49787 30251 49793
rect 30460 49827 30518 49833
rect 30460 49793 30472 49827
rect 30506 49824 30518 49827
rect 30926 49824 30932 49836
rect 30506 49796 30932 49824
rect 30506 49793 30518 49796
rect 30460 49787 30518 49793
rect 30926 49784 30932 49796
rect 30984 49784 30990 49836
rect 32030 49784 32036 49836
rect 32088 49824 32094 49836
rect 32125 49827 32183 49833
rect 32125 49824 32137 49827
rect 32088 49796 32137 49824
rect 32088 49784 32094 49796
rect 32125 49793 32137 49796
rect 32171 49793 32183 49827
rect 32125 49787 32183 49793
rect 32392 49827 32450 49833
rect 32392 49793 32404 49827
rect 32438 49824 32450 49827
rect 34238 49824 34244 49836
rect 32438 49796 34100 49824
rect 34199 49796 34244 49824
rect 32438 49793 32450 49796
rect 32392 49787 32450 49793
rect 29641 49759 29699 49765
rect 29641 49725 29653 49759
rect 29687 49756 29699 49759
rect 29730 49756 29736 49768
rect 29687 49728 29736 49756
rect 29687 49725 29699 49728
rect 29641 49719 29699 49725
rect 29730 49716 29736 49728
rect 29788 49716 29794 49768
rect 31386 49716 31392 49768
rect 31444 49756 31450 49768
rect 34072 49756 34100 49796
rect 34238 49784 34244 49796
rect 34296 49784 34302 49836
rect 35434 49824 35440 49836
rect 35395 49796 35440 49824
rect 35434 49784 35440 49796
rect 35492 49784 35498 49836
rect 35526 49784 35532 49836
rect 35584 49824 35590 49836
rect 35621 49827 35679 49833
rect 35621 49824 35633 49827
rect 35584 49796 35633 49824
rect 35584 49784 35590 49796
rect 35621 49793 35633 49796
rect 35667 49793 35679 49827
rect 35621 49787 35679 49793
rect 35713 49827 35771 49833
rect 35713 49793 35725 49827
rect 35759 49824 35771 49827
rect 35802 49824 35808 49836
rect 35759 49796 35808 49824
rect 35759 49793 35771 49796
rect 35713 49787 35771 49793
rect 35802 49784 35808 49796
rect 35860 49784 35866 49836
rect 36538 49824 36544 49836
rect 36499 49796 36544 49824
rect 36538 49784 36544 49796
rect 36596 49784 36602 49836
rect 37369 49827 37427 49833
rect 37369 49793 37381 49827
rect 37415 49793 37427 49827
rect 37476 49824 37504 49864
rect 37550 49852 37556 49904
rect 37608 49892 37614 49904
rect 38286 49892 38292 49904
rect 37608 49864 38292 49892
rect 37608 49852 37614 49864
rect 38286 49852 38292 49864
rect 38344 49852 38350 49904
rect 41690 49901 41696 49904
rect 41676 49895 41696 49901
rect 41676 49892 41688 49895
rect 38488 49864 39804 49892
rect 38488 49833 38516 49864
rect 38473 49827 38531 49833
rect 38473 49824 38485 49827
rect 37476 49796 38485 49824
rect 37369 49787 37427 49793
rect 38473 49793 38485 49796
rect 38519 49793 38531 49827
rect 38473 49787 38531 49793
rect 39485 49827 39543 49833
rect 39485 49793 39497 49827
rect 39531 49824 39543 49827
rect 39666 49824 39672 49836
rect 39531 49796 39672 49824
rect 39531 49793 39543 49796
rect 39485 49787 39543 49793
rect 36446 49756 36452 49768
rect 31444 49728 31616 49756
rect 34072 49728 36452 49756
rect 31444 49716 31450 49728
rect 31588 49697 31616 49728
rect 36446 49716 36452 49728
rect 36504 49716 36510 49768
rect 37090 49716 37096 49768
rect 37148 49756 37154 49768
rect 37384 49756 37412 49787
rect 39666 49784 39672 49796
rect 39724 49784 39730 49836
rect 39776 49756 39804 49864
rect 39960 49864 41688 49892
rect 39960 49833 39988 49864
rect 41676 49861 41688 49864
rect 41676 49855 41696 49861
rect 41690 49852 41696 49855
rect 41748 49852 41754 49904
rect 41800 49892 41828 49932
rect 42260 49932 43729 49960
rect 42260 49892 42288 49932
rect 43717 49929 43729 49932
rect 43763 49929 43775 49963
rect 43717 49923 43775 49929
rect 45922 49920 45928 49972
rect 45980 49960 45986 49972
rect 45980 49932 46336 49960
rect 45980 49920 45986 49932
rect 43349 49895 43407 49901
rect 43349 49892 43361 49895
rect 41800 49864 42288 49892
rect 42352 49864 43361 49892
rect 39945 49827 40003 49833
rect 39945 49793 39957 49827
rect 39991 49793 40003 49827
rect 42352 49824 42380 49864
rect 43349 49861 43361 49864
rect 43395 49892 43407 49895
rect 43438 49892 43444 49904
rect 43395 49864 43444 49892
rect 43395 49861 43407 49864
rect 43349 49855 43407 49861
rect 43438 49852 43444 49864
rect 43496 49852 43502 49904
rect 43533 49895 43591 49901
rect 43533 49861 43545 49895
rect 43579 49892 43591 49895
rect 44634 49892 44640 49904
rect 43579 49864 44640 49892
rect 43579 49861 43591 49864
rect 43533 49855 43591 49861
rect 44634 49852 44640 49864
rect 44692 49852 44698 49904
rect 44821 49895 44879 49901
rect 44821 49861 44833 49895
rect 44867 49892 44879 49895
rect 46308 49892 46336 49932
rect 46382 49920 46388 49972
rect 46440 49960 46446 49972
rect 46477 49963 46535 49969
rect 46477 49960 46489 49963
rect 46440 49932 46489 49960
rect 46440 49920 46446 49932
rect 46477 49929 46489 49932
rect 46523 49929 46535 49963
rect 49145 49963 49203 49969
rect 49145 49960 49157 49963
rect 46477 49923 46535 49929
rect 47596 49932 49157 49960
rect 47596 49892 47624 49932
rect 49145 49929 49157 49932
rect 49191 49929 49203 49963
rect 49145 49923 49203 49929
rect 49326 49920 49332 49972
rect 49384 49960 49390 49972
rect 50525 49963 50583 49969
rect 50525 49960 50537 49963
rect 49384 49932 50537 49960
rect 49384 49920 49390 49932
rect 50525 49929 50537 49932
rect 50571 49929 50583 49963
rect 51350 49960 51356 49972
rect 51311 49932 51356 49960
rect 50525 49923 50583 49929
rect 51350 49920 51356 49932
rect 51408 49920 51414 49972
rect 44867 49864 45968 49892
rect 46308 49864 47624 49892
rect 44867 49861 44879 49864
rect 44821 49855 44879 49861
rect 39945 49787 40003 49793
rect 40052 49822 41414 49824
rect 41524 49822 41644 49824
rect 41800 49822 42380 49824
rect 40052 49796 42380 49822
rect 40052 49756 40080 49796
rect 41386 49794 41552 49796
rect 41616 49794 41828 49796
rect 42426 49784 42432 49836
rect 42484 49824 42490 49836
rect 44729 49827 44787 49833
rect 42484 49796 42529 49824
rect 42484 49784 42490 49796
rect 44729 49793 44741 49827
rect 44775 49793 44787 49827
rect 44910 49824 44916 49836
rect 44871 49796 44916 49824
rect 44729 49787 44787 49793
rect 37148 49728 37412 49756
rect 38626 49728 39436 49756
rect 39776 49728 40080 49756
rect 40313 49759 40371 49765
rect 37148 49716 37154 49728
rect 31573 49691 31631 49697
rect 31573 49657 31585 49691
rect 31619 49657 31631 49691
rect 38626 49688 38654 49728
rect 39408 49697 39436 49728
rect 40313 49725 40325 49759
rect 40359 49756 40371 49759
rect 44545 49759 44603 49765
rect 44545 49756 44557 49759
rect 40359 49728 41644 49756
rect 40359 49725 40371 49728
rect 40313 49719 40371 49725
rect 31573 49651 31631 49657
rect 33051 49660 38654 49688
rect 39393 49691 39451 49697
rect 33051 49620 33079 49660
rect 39393 49657 39405 49691
rect 39439 49657 39451 49691
rect 41616 49688 41644 49728
rect 41800 49728 44557 49756
rect 41800 49688 41828 49728
rect 44545 49725 44557 49728
rect 44591 49725 44603 49759
rect 44545 49719 44603 49725
rect 39393 49651 39451 49657
rect 39500 49660 41460 49688
rect 41616 49660 41828 49688
rect 41877 49691 41935 49697
rect 29304 49592 33079 49620
rect 33502 49580 33508 49632
rect 33560 49620 33566 49632
rect 34609 49623 34667 49629
rect 34609 49620 34621 49623
rect 33560 49592 34621 49620
rect 33560 49580 33566 49592
rect 34609 49589 34621 49592
rect 34655 49589 34667 49623
rect 34790 49620 34796 49632
rect 34751 49592 34796 49620
rect 34609 49583 34667 49589
rect 34790 49580 34796 49592
rect 34848 49580 34854 49632
rect 37274 49580 37280 49632
rect 37332 49620 37338 49632
rect 39500 49620 39528 49660
rect 37332 49592 39528 49620
rect 41432 49620 41460 49660
rect 41877 49657 41889 49691
rect 41923 49688 41935 49691
rect 44174 49688 44180 49700
rect 41923 49660 44180 49688
rect 41923 49657 41935 49660
rect 41877 49651 41935 49657
rect 44174 49648 44180 49660
rect 44232 49648 44238 49700
rect 44744 49688 44772 49787
rect 44910 49784 44916 49796
rect 44968 49784 44974 49836
rect 45002 49784 45008 49836
rect 45060 49833 45066 49836
rect 45940 49833 45968 49864
rect 47670 49852 47676 49904
rect 47728 49892 47734 49904
rect 48133 49895 48191 49901
rect 48133 49892 48145 49895
rect 47728 49864 48145 49892
rect 47728 49852 47734 49864
rect 48133 49861 48145 49864
rect 48179 49892 48191 49895
rect 50065 49895 50123 49901
rect 50065 49892 50077 49895
rect 48179 49864 50077 49892
rect 48179 49861 48191 49864
rect 48133 49855 48191 49861
rect 50065 49861 50077 49864
rect 50111 49861 50123 49895
rect 50065 49855 50123 49861
rect 45060 49827 45089 49833
rect 45077 49793 45089 49827
rect 45060 49787 45089 49793
rect 45925 49827 45983 49833
rect 45925 49793 45937 49827
rect 45971 49824 45983 49827
rect 48777 49827 48835 49833
rect 45971 49796 48268 49824
rect 45971 49793 45983 49796
rect 45925 49787 45983 49793
rect 45060 49784 45066 49787
rect 45189 49759 45247 49765
rect 45189 49725 45201 49759
rect 45235 49756 45247 49759
rect 45646 49756 45652 49768
rect 45235 49728 45652 49756
rect 45235 49725 45247 49728
rect 45189 49719 45247 49725
rect 45646 49716 45652 49728
rect 45704 49716 45710 49768
rect 46201 49759 46259 49765
rect 46201 49725 46213 49759
rect 46247 49756 46259 49759
rect 46290 49756 46296 49768
rect 46247 49728 46296 49756
rect 46247 49725 46259 49728
rect 46201 49719 46259 49725
rect 46290 49716 46296 49728
rect 46348 49716 46354 49768
rect 47762 49756 47768 49768
rect 47723 49728 47768 49756
rect 47762 49716 47768 49728
rect 47820 49716 47826 49768
rect 45094 49688 45100 49700
rect 44744 49660 45100 49688
rect 45094 49648 45100 49660
rect 45152 49648 45158 49700
rect 48240 49688 48268 49796
rect 48777 49793 48789 49827
rect 48823 49824 48835 49827
rect 49326 49824 49332 49836
rect 48823 49796 49332 49824
rect 48823 49793 48835 49796
rect 48777 49787 48835 49793
rect 49326 49784 49332 49796
rect 49384 49784 49390 49836
rect 50341 49827 50399 49833
rect 50341 49793 50353 49827
rect 50387 49824 50399 49827
rect 50614 49824 50620 49836
rect 50387 49796 50620 49824
rect 50387 49793 50399 49796
rect 50341 49787 50399 49793
rect 50614 49784 50620 49796
rect 50672 49784 50678 49836
rect 51261 49827 51319 49833
rect 51261 49793 51273 49827
rect 51307 49824 51319 49827
rect 51350 49824 51356 49836
rect 51307 49796 51356 49824
rect 51307 49793 51319 49796
rect 51261 49787 51319 49793
rect 51350 49784 51356 49796
rect 51408 49784 51414 49836
rect 52086 49824 52092 49836
rect 52047 49796 52092 49824
rect 52086 49784 52092 49796
rect 52144 49784 52150 49836
rect 48869 49759 48927 49765
rect 48869 49756 48881 49759
rect 48424 49728 48881 49756
rect 48317 49691 48375 49697
rect 48317 49688 48329 49691
rect 48240 49660 48329 49688
rect 48317 49657 48329 49660
rect 48363 49657 48375 49691
rect 48317 49651 48375 49657
rect 42058 49620 42064 49632
rect 41432 49592 42064 49620
rect 37332 49580 37338 49592
rect 42058 49580 42064 49592
rect 42116 49580 42122 49632
rect 42610 49620 42616 49632
rect 42571 49592 42616 49620
rect 42610 49580 42616 49592
rect 42668 49580 42674 49632
rect 43530 49620 43536 49632
rect 43491 49592 43536 49620
rect 43530 49580 43536 49592
rect 43588 49580 43594 49632
rect 44910 49580 44916 49632
rect 44968 49620 44974 49632
rect 45370 49620 45376 49632
rect 44968 49592 45376 49620
rect 44968 49580 44974 49592
rect 45370 49580 45376 49592
rect 45428 49620 45434 49632
rect 46293 49623 46351 49629
rect 46293 49620 46305 49623
rect 45428 49592 46305 49620
rect 45428 49580 45434 49592
rect 46293 49589 46305 49592
rect 46339 49620 46351 49623
rect 46474 49620 46480 49632
rect 46339 49592 46480 49620
rect 46339 49589 46351 49592
rect 46293 49583 46351 49589
rect 46474 49580 46480 49592
rect 46532 49580 46538 49632
rect 48133 49623 48191 49629
rect 48133 49589 48145 49623
rect 48179 49620 48191 49623
rect 48222 49620 48228 49632
rect 48179 49592 48228 49620
rect 48179 49589 48191 49592
rect 48133 49583 48191 49589
rect 48222 49580 48228 49592
rect 48280 49620 48286 49632
rect 48424 49620 48452 49728
rect 48869 49725 48881 49728
rect 48915 49725 48927 49759
rect 50246 49756 50252 49768
rect 50207 49728 50252 49756
rect 48869 49719 48927 49725
rect 50246 49716 50252 49728
rect 50304 49716 50310 49768
rect 48280 49592 48452 49620
rect 48961 49623 49019 49629
rect 48280 49580 48286 49592
rect 48961 49589 48973 49623
rect 49007 49620 49019 49623
rect 49050 49620 49056 49632
rect 49007 49592 49056 49620
rect 49007 49589 49019 49592
rect 48961 49583 49019 49589
rect 49050 49580 49056 49592
rect 49108 49580 49114 49632
rect 50062 49620 50068 49632
rect 50023 49592 50068 49620
rect 50062 49580 50068 49592
rect 50120 49580 50126 49632
rect 51905 49623 51963 49629
rect 51905 49589 51917 49623
rect 51951 49620 51963 49623
rect 51994 49620 52000 49632
rect 51951 49592 52000 49620
rect 51951 49589 51963 49592
rect 51905 49583 51963 49589
rect 51994 49580 52000 49592
rect 52052 49580 52058 49632
rect 1104 49530 68816 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 65654 49530
rect 65706 49478 65718 49530
rect 65770 49478 65782 49530
rect 65834 49478 65846 49530
rect 65898 49478 65910 49530
rect 65962 49478 68816 49530
rect 1104 49456 68816 49478
rect 14366 49416 14372 49428
rect 14327 49388 14372 49416
rect 14366 49376 14372 49388
rect 14424 49376 14430 49428
rect 17586 49376 17592 49428
rect 17644 49416 17650 49428
rect 17681 49419 17739 49425
rect 17681 49416 17693 49419
rect 17644 49388 17693 49416
rect 17644 49376 17650 49388
rect 17681 49385 17693 49388
rect 17727 49385 17739 49419
rect 18506 49416 18512 49428
rect 18467 49388 18512 49416
rect 17681 49379 17739 49385
rect 13081 49283 13139 49289
rect 13081 49249 13093 49283
rect 13127 49280 13139 49283
rect 13814 49280 13820 49292
rect 13127 49252 13820 49280
rect 13127 49249 13139 49252
rect 13081 49243 13139 49249
rect 13814 49240 13820 49252
rect 13872 49240 13878 49292
rect 15378 49280 15384 49292
rect 14568 49252 15384 49280
rect 13262 49212 13268 49224
rect 13223 49184 13268 49212
rect 13262 49172 13268 49184
rect 13320 49172 13326 49224
rect 14568 49221 14596 49252
rect 15378 49240 15384 49252
rect 15436 49240 15442 49292
rect 17696 49280 17724 49379
rect 18506 49376 18512 49388
rect 18564 49376 18570 49428
rect 19334 49416 19340 49428
rect 19295 49388 19340 49416
rect 19334 49376 19340 49388
rect 19392 49376 19398 49428
rect 23014 49416 23020 49428
rect 22975 49388 23020 49416
rect 23014 49376 23020 49388
rect 23072 49376 23078 49428
rect 30926 49376 30932 49428
rect 30984 49416 30990 49428
rect 31113 49419 31171 49425
rect 31113 49416 31125 49419
rect 30984 49388 31125 49416
rect 30984 49376 30990 49388
rect 31113 49385 31125 49388
rect 31159 49385 31171 49419
rect 31113 49379 31171 49385
rect 31220 49388 31754 49416
rect 28718 49308 28724 49360
rect 28776 49348 28782 49360
rect 31220 49348 31248 49388
rect 28776 49320 31248 49348
rect 28776 49308 28782 49320
rect 18141 49283 18199 49289
rect 18141 49280 18153 49283
rect 17696 49252 18153 49280
rect 18141 49249 18153 49252
rect 18187 49249 18199 49283
rect 20165 49283 20223 49289
rect 20165 49280 20177 49283
rect 18141 49243 18199 49249
rect 18340 49252 20177 49280
rect 14553 49215 14611 49221
rect 14553 49181 14565 49215
rect 14599 49181 14611 49215
rect 14553 49175 14611 49181
rect 15013 49215 15071 49221
rect 15013 49181 15025 49215
rect 15059 49181 15071 49215
rect 15013 49175 15071 49181
rect 15028 49144 15056 49175
rect 15194 49172 15200 49224
rect 15252 49212 15258 49224
rect 15289 49215 15347 49221
rect 15289 49212 15301 49215
rect 15252 49184 15301 49212
rect 15252 49172 15258 49184
rect 15289 49181 15301 49184
rect 15335 49181 15347 49215
rect 15289 49175 15347 49181
rect 16301 49215 16359 49221
rect 16301 49181 16313 49215
rect 16347 49212 16359 49215
rect 16850 49212 16856 49224
rect 16347 49184 16856 49212
rect 16347 49181 16359 49184
rect 16301 49175 16359 49181
rect 16850 49172 16856 49184
rect 16908 49172 16914 49224
rect 17310 49172 17316 49224
rect 17368 49212 17374 49224
rect 18340 49221 18368 49252
rect 20165 49249 20177 49252
rect 20211 49249 20223 49283
rect 31726 49280 31754 49388
rect 35434 49376 35440 49428
rect 35492 49416 35498 49428
rect 36081 49419 36139 49425
rect 36081 49416 36093 49419
rect 35492 49388 36093 49416
rect 35492 49376 35498 49388
rect 36081 49385 36093 49388
rect 36127 49385 36139 49419
rect 36081 49379 36139 49385
rect 39117 49419 39175 49425
rect 39117 49385 39129 49419
rect 39163 49416 39175 49419
rect 40034 49416 40040 49428
rect 39163 49388 40040 49416
rect 39163 49385 39175 49388
rect 39117 49379 39175 49385
rect 40034 49376 40040 49388
rect 40092 49416 40098 49428
rect 41322 49416 41328 49428
rect 40092 49388 41328 49416
rect 40092 49376 40098 49388
rect 41322 49376 41328 49388
rect 41380 49376 41386 49428
rect 43530 49376 43536 49428
rect 43588 49416 43594 49428
rect 46290 49416 46296 49428
rect 43588 49388 46152 49416
rect 46251 49388 46296 49416
rect 43588 49376 43594 49388
rect 40126 49348 40132 49360
rect 35728 49320 39988 49348
rect 40087 49320 40132 49348
rect 31726 49252 34836 49280
rect 20165 49243 20223 49249
rect 18325 49215 18383 49221
rect 18325 49212 18337 49215
rect 17368 49184 18337 49212
rect 17368 49172 17374 49184
rect 18325 49181 18337 49184
rect 18371 49181 18383 49215
rect 18325 49175 18383 49181
rect 19245 49215 19303 49221
rect 19245 49181 19257 49215
rect 19291 49181 19303 49215
rect 19245 49175 19303 49181
rect 19889 49215 19947 49221
rect 19889 49181 19901 49215
rect 19935 49212 19947 49215
rect 20530 49212 20536 49224
rect 19935 49184 20536 49212
rect 19935 49181 19947 49184
rect 19889 49175 19947 49181
rect 16022 49144 16028 49156
rect 15028 49116 16028 49144
rect 16022 49104 16028 49116
rect 16080 49104 16086 49156
rect 16574 49153 16580 49156
rect 16568 49107 16580 49153
rect 16632 49144 16638 49156
rect 19260 49144 19288 49175
rect 20530 49172 20536 49184
rect 20588 49172 20594 49224
rect 21637 49215 21695 49221
rect 21637 49181 21649 49215
rect 21683 49212 21695 49215
rect 22186 49212 22192 49224
rect 21683 49184 22192 49212
rect 21683 49181 21695 49184
rect 21637 49175 21695 49181
rect 22186 49172 22192 49184
rect 22244 49172 22250 49224
rect 23290 49172 23296 49224
rect 23348 49172 23354 49224
rect 24854 49212 24860 49224
rect 24815 49184 24860 49212
rect 24854 49172 24860 49184
rect 24912 49172 24918 49224
rect 24949 49215 25007 49221
rect 24949 49181 24961 49215
rect 24995 49212 25007 49215
rect 25501 49215 25559 49221
rect 25501 49212 25513 49215
rect 24995 49184 25513 49212
rect 24995 49181 25007 49184
rect 24949 49175 25007 49181
rect 25501 49181 25513 49184
rect 25547 49181 25559 49215
rect 25501 49175 25559 49181
rect 25768 49215 25826 49221
rect 25768 49181 25780 49215
rect 25814 49212 25826 49215
rect 26050 49212 26056 49224
rect 25814 49184 26056 49212
rect 25814 49181 25826 49184
rect 25768 49175 25826 49181
rect 26050 49172 26056 49184
rect 26108 49172 26114 49224
rect 26326 49172 26332 49224
rect 26384 49212 26390 49224
rect 27617 49215 27675 49221
rect 27617 49212 27629 49215
rect 26384 49184 27629 49212
rect 26384 49172 26390 49184
rect 27617 49181 27629 49184
rect 27663 49181 27675 49215
rect 27617 49175 27675 49181
rect 27884 49215 27942 49221
rect 27884 49181 27896 49215
rect 27930 49212 27942 49215
rect 28626 49212 28632 49224
rect 27930 49184 28632 49212
rect 27930 49181 27942 49184
rect 27884 49175 27942 49181
rect 28626 49172 28632 49184
rect 28684 49172 28690 49224
rect 30282 49212 30288 49224
rect 30243 49184 30288 49212
rect 30282 49172 30288 49184
rect 30340 49172 30346 49224
rect 31294 49212 31300 49224
rect 31255 49184 31300 49212
rect 31294 49172 31300 49184
rect 31352 49172 31358 49224
rect 32582 49212 32588 49224
rect 32543 49184 32588 49212
rect 32582 49172 32588 49184
rect 32640 49172 32646 49224
rect 34698 49212 34704 49224
rect 34659 49184 34704 49212
rect 34698 49172 34704 49184
rect 34756 49172 34762 49224
rect 34808 49212 34836 49252
rect 35728 49212 35756 49320
rect 38381 49283 38439 49289
rect 38381 49249 38393 49283
rect 38427 49280 38439 49283
rect 38427 49252 39712 49280
rect 38427 49249 38439 49252
rect 38381 49243 38439 49249
rect 39684 49224 39712 49252
rect 34808 49184 35756 49212
rect 36630 49172 36636 49224
rect 36688 49212 36694 49224
rect 37093 49215 37151 49221
rect 37093 49212 37105 49215
rect 36688 49184 37105 49212
rect 36688 49172 36694 49184
rect 37093 49181 37105 49184
rect 37139 49212 37151 49215
rect 37139 49184 38240 49212
rect 37139 49181 37151 49184
rect 37093 49175 37151 49181
rect 20254 49144 20260 49156
rect 16632 49116 16668 49144
rect 19260 49116 20260 49144
rect 16574 49104 16580 49107
rect 16632 49104 16638 49116
rect 20254 49104 20260 49116
rect 20312 49104 20318 49156
rect 21904 49147 21962 49153
rect 21904 49113 21916 49147
rect 21950 49144 21962 49147
rect 22370 49144 22376 49156
rect 21950 49116 22376 49144
rect 21950 49113 21962 49116
rect 21904 49107 21962 49113
rect 22370 49104 22376 49116
rect 22428 49104 22434 49156
rect 23308 49144 23336 49172
rect 30653 49147 30711 49153
rect 30653 49144 30665 49147
rect 23308 49116 30665 49144
rect 30653 49113 30665 49116
rect 30699 49144 30711 49147
rect 30834 49144 30840 49156
rect 30699 49116 30840 49144
rect 30699 49113 30711 49116
rect 30653 49107 30711 49113
rect 30834 49104 30840 49116
rect 30892 49104 30898 49156
rect 32674 49104 32680 49156
rect 32732 49144 32738 49156
rect 32953 49147 33011 49153
rect 32953 49144 32965 49147
rect 32732 49116 32965 49144
rect 32732 49104 32738 49116
rect 32953 49113 32965 49116
rect 32999 49144 33011 49147
rect 33042 49144 33048 49156
rect 32999 49116 33048 49144
rect 32999 49113 33011 49116
rect 32953 49107 33011 49113
rect 33042 49104 33048 49116
rect 33100 49104 33106 49156
rect 33410 49104 33416 49156
rect 33468 49144 33474 49156
rect 33597 49147 33655 49153
rect 33597 49144 33609 49147
rect 33468 49116 33609 49144
rect 33468 49104 33474 49116
rect 33597 49113 33609 49116
rect 33643 49113 33655 49147
rect 33597 49107 33655 49113
rect 34606 49104 34612 49156
rect 34664 49144 34670 49156
rect 34946 49147 35004 49153
rect 34946 49144 34958 49147
rect 34664 49116 34958 49144
rect 34664 49104 34670 49116
rect 34946 49113 34958 49116
rect 34992 49113 35004 49147
rect 34946 49107 35004 49113
rect 36538 49104 36544 49156
rect 36596 49144 36602 49156
rect 37642 49144 37648 49156
rect 36596 49116 37648 49144
rect 36596 49104 36602 49116
rect 37642 49104 37648 49116
rect 37700 49104 37706 49156
rect 13170 49036 13176 49088
rect 13228 49076 13234 49088
rect 13449 49079 13507 49085
rect 13449 49076 13461 49079
rect 13228 49048 13461 49076
rect 13228 49036 13234 49048
rect 13449 49045 13461 49048
rect 13495 49045 13507 49079
rect 16040 49076 16068 49104
rect 23290 49076 23296 49088
rect 16040 49048 23296 49076
rect 13449 49039 13507 49045
rect 23290 49036 23296 49048
rect 23348 49036 23354 49088
rect 26881 49079 26939 49085
rect 26881 49045 26893 49079
rect 26927 49076 26939 49079
rect 27614 49076 27620 49088
rect 26927 49048 27620 49076
rect 26927 49045 26939 49048
rect 26881 49039 26939 49045
rect 27614 49036 27620 49048
rect 27672 49036 27678 49088
rect 28997 49079 29055 49085
rect 28997 49045 29009 49079
rect 29043 49076 29055 49079
rect 29086 49076 29092 49088
rect 29043 49048 29092 49076
rect 29043 49045 29055 49048
rect 28997 49039 29055 49045
rect 29086 49036 29092 49048
rect 29144 49036 29150 49088
rect 33502 49036 33508 49088
rect 33560 49076 33566 49088
rect 33689 49079 33747 49085
rect 33689 49076 33701 49079
rect 33560 49048 33701 49076
rect 33560 49036 33566 49048
rect 33689 49045 33701 49048
rect 33735 49045 33747 49079
rect 37274 49076 37280 49088
rect 37187 49048 37280 49076
rect 33689 49039 33747 49045
rect 37274 49036 37280 49048
rect 37332 49076 37338 49088
rect 37458 49076 37464 49088
rect 37332 49048 37464 49076
rect 37332 49036 37338 49048
rect 37458 49036 37464 49048
rect 37516 49036 37522 49088
rect 38212 49076 38240 49184
rect 38286 49172 38292 49224
rect 38344 49212 38350 49224
rect 38933 49215 38991 49221
rect 38344 49184 38389 49212
rect 38344 49172 38350 49184
rect 38933 49181 38945 49215
rect 38979 49181 38991 49215
rect 38933 49175 38991 49181
rect 38948 49076 38976 49175
rect 39666 49172 39672 49224
rect 39724 49212 39730 49224
rect 39853 49215 39911 49221
rect 39853 49212 39865 49215
rect 39724 49184 39865 49212
rect 39724 49172 39730 49184
rect 39853 49181 39865 49184
rect 39899 49181 39911 49215
rect 39853 49175 39911 49181
rect 39960 49144 39988 49320
rect 40126 49308 40132 49320
rect 40184 49308 40190 49360
rect 41690 49348 41696 49360
rect 40788 49320 41696 49348
rect 40589 49215 40647 49221
rect 40589 49181 40601 49215
rect 40635 49212 40647 49215
rect 40788 49212 40816 49320
rect 41690 49308 41696 49320
rect 41748 49348 41754 49360
rect 42610 49348 42616 49360
rect 41748 49320 42616 49348
rect 41748 49308 41754 49320
rect 42610 49308 42616 49320
rect 42668 49308 42674 49360
rect 45554 49348 45560 49360
rect 43732 49320 45560 49348
rect 40865 49283 40923 49289
rect 40865 49249 40877 49283
rect 40911 49280 40923 49283
rect 40911 49252 43208 49280
rect 40911 49249 40923 49252
rect 40865 49243 40923 49249
rect 40635 49184 40816 49212
rect 40635 49181 40647 49184
rect 40589 49175 40647 49181
rect 41414 49172 41420 49224
rect 41472 49212 41478 49224
rect 41601 49215 41659 49221
rect 41472 49184 41517 49212
rect 41472 49172 41478 49184
rect 41601 49181 41613 49215
rect 41647 49212 41659 49215
rect 41690 49212 41696 49224
rect 41647 49184 41696 49212
rect 41647 49181 41659 49184
rect 41601 49175 41659 49181
rect 41690 49172 41696 49184
rect 41748 49172 41754 49224
rect 41966 49212 41972 49224
rect 41927 49184 41972 49212
rect 41966 49172 41972 49184
rect 42024 49172 42030 49224
rect 42889 49147 42947 49153
rect 42889 49144 42901 49147
rect 39960 49116 42901 49144
rect 42889 49113 42901 49116
rect 42935 49113 42947 49147
rect 43180 49144 43208 49252
rect 43438 49212 43444 49224
rect 43399 49184 43444 49212
rect 43438 49172 43444 49184
rect 43496 49172 43502 49224
rect 43732 49221 43760 49320
rect 45554 49308 45560 49320
rect 45612 49308 45618 49360
rect 46124 49348 46152 49388
rect 46290 49376 46296 49388
rect 46348 49376 46354 49428
rect 48314 49376 48320 49428
rect 48372 49416 48378 49428
rect 48777 49419 48835 49425
rect 48777 49416 48789 49419
rect 48372 49388 48789 49416
rect 48372 49376 48378 49388
rect 48777 49385 48789 49388
rect 48823 49385 48835 49419
rect 48777 49379 48835 49385
rect 51261 49419 51319 49425
rect 51261 49385 51273 49419
rect 51307 49416 51319 49419
rect 52086 49416 52092 49428
rect 51307 49388 52092 49416
rect 51307 49385 51319 49388
rect 51261 49379 51319 49385
rect 52086 49376 52092 49388
rect 52144 49376 52150 49428
rect 47486 49348 47492 49360
rect 46124 49320 47492 49348
rect 47486 49308 47492 49320
rect 47544 49308 47550 49360
rect 45204 49252 46152 49280
rect 43717 49215 43775 49221
rect 43717 49181 43729 49215
rect 43763 49181 43775 49215
rect 43898 49212 43904 49224
rect 43859 49184 43904 49212
rect 43717 49175 43775 49181
rect 43898 49172 43904 49184
rect 43956 49172 43962 49224
rect 45204 49221 45232 49252
rect 45189 49215 45247 49221
rect 45189 49181 45201 49215
rect 45235 49181 45247 49215
rect 45370 49212 45376 49224
rect 45331 49184 45376 49212
rect 45189 49175 45247 49181
rect 45370 49172 45376 49184
rect 45428 49172 45434 49224
rect 45646 49212 45652 49224
rect 45607 49184 45652 49212
rect 45646 49172 45652 49184
rect 45704 49172 45710 49224
rect 46124 49221 46152 49252
rect 48700 49252 49556 49280
rect 46109 49215 46167 49221
rect 46109 49181 46121 49215
rect 46155 49181 46167 49215
rect 46474 49212 46480 49224
rect 46387 49184 46480 49212
rect 46109 49175 46167 49181
rect 45005 49147 45063 49153
rect 45005 49144 45017 49147
rect 43180 49116 45017 49144
rect 42889 49107 42947 49113
rect 45005 49113 45017 49116
rect 45051 49113 45063 49147
rect 45005 49107 45063 49113
rect 45094 49104 45100 49156
rect 45152 49144 45158 49156
rect 45281 49147 45339 49153
rect 45281 49144 45293 49147
rect 45152 49116 45293 49144
rect 45152 49104 45158 49116
rect 45281 49113 45293 49116
rect 45327 49113 45339 49147
rect 45281 49107 45339 49113
rect 45491 49147 45549 49153
rect 45491 49113 45503 49147
rect 45537 49113 45549 49147
rect 46124 49144 46152 49175
rect 46474 49172 46480 49184
rect 46532 49212 46538 49224
rect 47670 49212 47676 49224
rect 46532 49184 47676 49212
rect 46532 49172 46538 49184
rect 47670 49172 47676 49184
rect 47728 49172 47734 49224
rect 48590 49172 48596 49224
rect 48648 49212 48654 49224
rect 48700 49221 48728 49252
rect 48685 49215 48743 49221
rect 48685 49212 48697 49215
rect 48648 49184 48697 49212
rect 48648 49172 48654 49184
rect 48685 49181 48697 49184
rect 48731 49181 48743 49215
rect 49326 49212 49332 49224
rect 49287 49184 49332 49212
rect 48685 49175 48743 49181
rect 49326 49172 49332 49184
rect 49384 49172 49390 49224
rect 49528 49221 49556 49252
rect 49513 49215 49571 49221
rect 49513 49181 49525 49215
rect 49559 49181 49571 49215
rect 49513 49175 49571 49181
rect 50246 49172 50252 49224
rect 50304 49212 50310 49224
rect 50985 49215 51043 49221
rect 50985 49212 50997 49215
rect 50304 49184 50997 49212
rect 50304 49172 50310 49184
rect 50985 49181 50997 49184
rect 51031 49181 51043 49215
rect 50985 49175 51043 49181
rect 51077 49215 51135 49221
rect 51077 49181 51089 49215
rect 51123 49212 51135 49215
rect 51534 49212 51540 49224
rect 51123 49184 51540 49212
rect 51123 49181 51135 49184
rect 51077 49175 51135 49181
rect 49421 49147 49479 49153
rect 49421 49144 49433 49147
rect 46124 49116 49433 49144
rect 45491 49107 45549 49113
rect 49421 49113 49433 49116
rect 49467 49113 49479 49147
rect 49421 49107 49479 49113
rect 40218 49076 40224 49088
rect 38212 49048 40224 49076
rect 40218 49036 40224 49048
rect 40276 49036 40282 49088
rect 40310 49036 40316 49088
rect 40368 49076 40374 49088
rect 41601 49079 41659 49085
rect 41601 49076 41613 49079
rect 40368 49048 41613 49076
rect 40368 49036 40374 49048
rect 41601 49045 41613 49048
rect 41647 49045 41659 49079
rect 41601 49039 41659 49045
rect 45370 49036 45376 49088
rect 45428 49076 45434 49088
rect 45506 49076 45534 49107
rect 45428 49048 45534 49076
rect 45428 49036 45434 49048
rect 45922 49036 45928 49088
rect 45980 49076 45986 49088
rect 46661 49079 46719 49085
rect 46661 49076 46673 49079
rect 45980 49048 46673 49076
rect 45980 49036 45986 49048
rect 46661 49045 46673 49048
rect 46707 49045 46719 49079
rect 51000 49076 51028 49175
rect 51534 49172 51540 49184
rect 51592 49172 51598 49224
rect 51626 49172 51632 49224
rect 51684 49212 51690 49224
rect 51994 49221 52000 49224
rect 51721 49215 51779 49221
rect 51721 49212 51733 49215
rect 51684 49184 51733 49212
rect 51684 49172 51690 49184
rect 51721 49181 51733 49184
rect 51767 49181 51779 49215
rect 51988 49212 52000 49221
rect 51955 49184 52000 49212
rect 51721 49175 51779 49181
rect 51988 49175 52000 49184
rect 51994 49172 52000 49175
rect 52052 49172 52058 49224
rect 53101 49079 53159 49085
rect 53101 49076 53113 49079
rect 51000 49048 53113 49076
rect 46661 49039 46719 49045
rect 53101 49045 53113 49048
rect 53147 49045 53159 49079
rect 53101 49039 53159 49045
rect 1104 48986 68816 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 68816 48986
rect 1104 48912 68816 48934
rect 12986 48872 12992 48884
rect 12947 48844 12992 48872
rect 12986 48832 12992 48844
rect 13044 48832 13050 48884
rect 19613 48875 19671 48881
rect 19613 48841 19625 48875
rect 19659 48872 19671 48875
rect 20714 48872 20720 48884
rect 19659 48844 20720 48872
rect 19659 48841 19671 48844
rect 19613 48835 19671 48841
rect 20714 48832 20720 48844
rect 20772 48832 20778 48884
rect 21177 48875 21235 48881
rect 21177 48841 21189 48875
rect 21223 48841 21235 48875
rect 26326 48872 26332 48884
rect 26287 48844 26332 48872
rect 21177 48835 21235 48841
rect 13262 48764 13268 48816
rect 13320 48804 13326 48816
rect 17313 48807 17371 48813
rect 17313 48804 17325 48807
rect 13320 48776 17325 48804
rect 13320 48764 13326 48776
rect 17313 48773 17325 48776
rect 17359 48773 17371 48807
rect 20806 48804 20812 48816
rect 17313 48767 17371 48773
rect 20272 48776 20812 48804
rect 20272 48748 20300 48776
rect 20806 48764 20812 48776
rect 20864 48804 20870 48816
rect 21192 48804 21220 48835
rect 26326 48832 26332 48844
rect 26384 48832 26390 48884
rect 27338 48872 27344 48884
rect 27299 48844 27344 48872
rect 27338 48832 27344 48844
rect 27396 48832 27402 48884
rect 29178 48832 29184 48884
rect 29236 48872 29242 48884
rect 29457 48875 29515 48881
rect 29457 48872 29469 48875
rect 29236 48844 29469 48872
rect 29236 48832 29242 48844
rect 29457 48841 29469 48844
rect 29503 48841 29515 48875
rect 34606 48872 34612 48884
rect 34567 48844 34612 48872
rect 29457 48835 29515 48841
rect 34606 48832 34612 48844
rect 34664 48832 34670 48884
rect 36541 48875 36599 48881
rect 36541 48841 36553 48875
rect 36587 48841 36599 48875
rect 41414 48872 41420 48884
rect 36541 48835 36599 48841
rect 27982 48804 27988 48816
rect 20864 48776 21220 48804
rect 24780 48776 27988 48804
rect 20864 48764 20870 48776
rect 13170 48736 13176 48748
rect 13131 48708 13176 48736
rect 13170 48696 13176 48708
rect 13228 48696 13234 48748
rect 14001 48739 14059 48745
rect 14001 48705 14013 48739
rect 14047 48736 14059 48739
rect 17126 48736 17132 48748
rect 14047 48708 16574 48736
rect 17087 48708 17132 48736
rect 14047 48705 14059 48708
rect 14001 48699 14059 48705
rect 16546 48600 16574 48708
rect 17126 48696 17132 48708
rect 17184 48696 17190 48748
rect 19797 48739 19855 48745
rect 19797 48705 19809 48739
rect 19843 48736 19855 48739
rect 19978 48736 19984 48748
rect 19843 48708 19984 48736
rect 19843 48705 19855 48708
rect 19797 48699 19855 48705
rect 19978 48696 19984 48708
rect 20036 48696 20042 48748
rect 20254 48736 20260 48748
rect 20215 48708 20260 48736
rect 20254 48696 20260 48708
rect 20312 48696 20318 48748
rect 20990 48736 20996 48748
rect 20951 48708 20996 48736
rect 20990 48696 20996 48708
rect 21048 48696 21054 48748
rect 24780 48745 24808 48776
rect 27982 48764 27988 48776
rect 28040 48764 28046 48816
rect 29086 48804 29092 48816
rect 29047 48776 29092 48804
rect 29086 48764 29092 48776
rect 29144 48764 29150 48816
rect 29289 48807 29347 48813
rect 29289 48804 29301 48807
rect 29288 48773 29301 48804
rect 29335 48804 29347 48807
rect 29546 48804 29552 48816
rect 29335 48776 29552 48804
rect 29335 48773 29347 48776
rect 29288 48767 29347 48773
rect 24765 48739 24823 48745
rect 24765 48736 24777 48739
rect 22848 48708 24777 48736
rect 20530 48628 20536 48680
rect 20588 48668 20594 48680
rect 22848 48668 22876 48708
rect 24765 48705 24777 48708
rect 24811 48705 24823 48739
rect 24765 48699 24823 48705
rect 24949 48739 25007 48745
rect 24949 48705 24961 48739
rect 24995 48736 25007 48739
rect 25593 48739 25651 48745
rect 25593 48736 25605 48739
rect 24995 48708 25605 48736
rect 24995 48705 25007 48708
rect 24949 48699 25007 48705
rect 25593 48705 25605 48708
rect 25639 48705 25651 48739
rect 25593 48699 25651 48705
rect 26237 48739 26295 48745
rect 26237 48705 26249 48739
rect 26283 48736 26295 48739
rect 26510 48736 26516 48748
rect 26283 48708 26516 48736
rect 26283 48705 26295 48708
rect 26237 48699 26295 48705
rect 26510 48696 26516 48708
rect 26568 48696 26574 48748
rect 27157 48739 27215 48745
rect 27157 48705 27169 48739
rect 27203 48736 27215 48739
rect 27890 48736 27896 48748
rect 27203 48708 27896 48736
rect 27203 48705 27215 48708
rect 27157 48699 27215 48705
rect 27890 48696 27896 48708
rect 27948 48736 27954 48748
rect 28718 48736 28724 48748
rect 27948 48708 28724 48736
rect 27948 48696 27954 48708
rect 28718 48696 28724 48708
rect 28776 48696 28782 48748
rect 28813 48739 28871 48745
rect 28813 48705 28825 48739
rect 28859 48736 28871 48739
rect 29288 48736 29316 48767
rect 29546 48764 29552 48776
rect 29604 48764 29610 48816
rect 30009 48807 30067 48813
rect 30009 48773 30021 48807
rect 30055 48804 30067 48807
rect 30282 48804 30288 48816
rect 30055 48776 30288 48804
rect 30055 48773 30067 48776
rect 30009 48767 30067 48773
rect 30282 48764 30288 48776
rect 30340 48764 30346 48816
rect 36556 48804 36584 48835
rect 41386 48832 41420 48872
rect 41472 48872 41478 48884
rect 41693 48875 41751 48881
rect 41693 48872 41705 48875
rect 41472 48844 41705 48872
rect 41472 48832 41478 48844
rect 41693 48841 41705 48844
rect 41739 48841 41751 48875
rect 41693 48835 41751 48841
rect 42610 48832 42616 48884
rect 42668 48872 42674 48884
rect 43898 48872 43904 48884
rect 42668 48844 43300 48872
rect 43859 48844 43904 48872
rect 42668 48832 42674 48844
rect 37522 48807 37580 48813
rect 37522 48804 37534 48807
rect 36556 48776 37534 48804
rect 37522 48773 37534 48776
rect 37568 48773 37580 48807
rect 41386 48804 41414 48832
rect 37522 48767 37580 48773
rect 39960 48776 41414 48804
rect 34790 48736 34796 48748
rect 28859 48708 29316 48736
rect 34751 48708 34796 48736
rect 28859 48705 28871 48708
rect 28813 48699 28871 48705
rect 34790 48696 34796 48708
rect 34848 48696 34854 48748
rect 36725 48739 36783 48745
rect 36725 48705 36737 48739
rect 36771 48736 36783 48739
rect 37366 48736 37372 48748
rect 36771 48708 37372 48736
rect 36771 48705 36783 48708
rect 36725 48699 36783 48705
rect 37366 48696 37372 48708
rect 37424 48696 37430 48748
rect 39960 48745 39988 48776
rect 43162 48764 43168 48816
rect 43220 48764 43226 48816
rect 43272 48804 43300 48844
rect 43898 48832 43904 48844
rect 43956 48832 43962 48884
rect 45922 48872 45928 48884
rect 45883 48844 45928 48872
rect 45922 48832 45928 48844
rect 45980 48832 45986 48884
rect 46014 48832 46020 48884
rect 46072 48872 46078 48884
rect 46934 48872 46940 48884
rect 46072 48844 46117 48872
rect 46895 48844 46940 48872
rect 46072 48832 46078 48844
rect 46934 48832 46940 48844
rect 46992 48832 46998 48884
rect 47791 48875 47849 48881
rect 47791 48872 47803 48875
rect 47044 48844 47803 48872
rect 43272 48776 43944 48804
rect 39853 48739 39911 48745
rect 39853 48705 39865 48739
rect 39899 48705 39911 48739
rect 39853 48699 39911 48705
rect 39945 48739 40003 48745
rect 39945 48705 39957 48739
rect 39991 48705 40003 48739
rect 39945 48699 40003 48705
rect 40681 48739 40739 48745
rect 40681 48705 40693 48739
rect 40727 48736 40739 48739
rect 41509 48739 41567 48745
rect 40727 48708 41460 48736
rect 40727 48705 40739 48708
rect 40681 48699 40739 48705
rect 20588 48640 22876 48668
rect 24581 48671 24639 48677
rect 20588 48628 20594 48640
rect 24581 48637 24593 48671
rect 24627 48668 24639 48671
rect 24854 48668 24860 48680
rect 24627 48640 24860 48668
rect 24627 48637 24639 48640
rect 24581 48631 24639 48637
rect 24854 48628 24860 48640
rect 24912 48628 24918 48680
rect 26973 48671 27031 48677
rect 26973 48637 26985 48671
rect 27019 48668 27031 48671
rect 27614 48668 27620 48680
rect 27019 48640 27620 48668
rect 27019 48637 27031 48640
rect 26973 48631 27031 48637
rect 27614 48628 27620 48640
rect 27672 48668 27678 48680
rect 28442 48668 28448 48680
rect 27672 48640 28448 48668
rect 27672 48628 27678 48640
rect 28442 48628 28448 48640
rect 28500 48628 28506 48680
rect 34698 48628 34704 48680
rect 34756 48668 34762 48680
rect 37277 48671 37335 48677
rect 37277 48668 37289 48671
rect 34756 48640 37289 48668
rect 34756 48628 34762 48640
rect 37277 48637 37289 48640
rect 37323 48637 37335 48671
rect 37277 48631 37335 48637
rect 30098 48600 30104 48612
rect 16546 48572 30104 48600
rect 30098 48560 30104 48572
rect 30156 48600 30162 48612
rect 30193 48603 30251 48609
rect 30193 48600 30205 48603
rect 30156 48572 30205 48600
rect 30156 48560 30162 48572
rect 30193 48569 30205 48572
rect 30239 48569 30251 48603
rect 30193 48563 30251 48569
rect 14090 48492 14096 48544
rect 14148 48532 14154 48544
rect 14185 48535 14243 48541
rect 14185 48532 14197 48535
rect 14148 48504 14197 48532
rect 14148 48492 14154 48504
rect 14185 48501 14197 48504
rect 14231 48501 14243 48535
rect 20438 48532 20444 48544
rect 20399 48504 20444 48532
rect 14185 48495 14243 48501
rect 20438 48492 20444 48504
rect 20496 48492 20502 48544
rect 25406 48532 25412 48544
rect 25367 48504 25412 48532
rect 25406 48492 25412 48504
rect 25464 48492 25470 48544
rect 29273 48535 29331 48541
rect 29273 48501 29285 48535
rect 29319 48532 29331 48535
rect 30006 48532 30012 48544
rect 29319 48504 30012 48532
rect 29319 48501 29331 48504
rect 29273 48495 29331 48501
rect 30006 48492 30012 48504
rect 30064 48492 30070 48544
rect 33410 48492 33416 48544
rect 33468 48532 33474 48544
rect 37550 48532 37556 48544
rect 33468 48504 37556 48532
rect 33468 48492 33474 48504
rect 37550 48492 37556 48504
rect 37608 48492 37614 48544
rect 37918 48492 37924 48544
rect 37976 48532 37982 48544
rect 38657 48535 38715 48541
rect 38657 48532 38669 48535
rect 37976 48504 38669 48532
rect 37976 48492 37982 48504
rect 38657 48501 38669 48504
rect 38703 48501 38715 48535
rect 39868 48532 39896 48699
rect 40129 48671 40187 48677
rect 40129 48637 40141 48671
rect 40175 48668 40187 48671
rect 40218 48668 40224 48680
rect 40175 48640 40224 48668
rect 40175 48637 40187 48640
rect 40129 48631 40187 48637
rect 40218 48628 40224 48640
rect 40276 48628 40282 48680
rect 41322 48668 41328 48680
rect 41283 48640 41328 48668
rect 41322 48628 41328 48640
rect 41380 48628 41386 48680
rect 41432 48668 41460 48708
rect 41509 48705 41521 48739
rect 41555 48736 41567 48739
rect 41598 48736 41604 48748
rect 41555 48708 41604 48736
rect 41555 48705 41567 48708
rect 41509 48699 41567 48705
rect 41598 48696 41604 48708
rect 41656 48736 41662 48748
rect 42978 48736 42984 48748
rect 41656 48708 42840 48736
rect 42939 48708 42984 48736
rect 41656 48696 41662 48708
rect 41782 48668 41788 48680
rect 41432 48640 41788 48668
rect 41782 48628 41788 48640
rect 41840 48628 41846 48680
rect 42812 48677 42840 48708
rect 42978 48696 42984 48708
rect 43036 48696 43042 48748
rect 42797 48671 42855 48677
rect 42797 48637 42809 48671
rect 42843 48637 42855 48671
rect 43070 48668 43076 48680
rect 43031 48640 43076 48668
rect 42797 48631 42855 48637
rect 43070 48628 43076 48640
rect 43128 48628 43134 48680
rect 43180 48677 43208 48764
rect 43714 48736 43720 48748
rect 43675 48708 43720 48736
rect 43714 48696 43720 48708
rect 43772 48696 43778 48748
rect 43916 48745 43944 48776
rect 45738 48764 45744 48816
rect 45796 48804 45802 48816
rect 45833 48807 45891 48813
rect 45833 48804 45845 48807
rect 45796 48776 45845 48804
rect 45796 48764 45802 48776
rect 45833 48773 45845 48776
rect 45879 48773 45891 48807
rect 47044 48804 47072 48844
rect 47791 48841 47803 48844
rect 47837 48872 47849 48875
rect 48130 48872 48136 48884
rect 47837 48844 48136 48872
rect 47837 48841 47849 48844
rect 47791 48835 47849 48841
rect 48130 48832 48136 48844
rect 48188 48832 48194 48884
rect 51626 48872 51632 48884
rect 51587 48844 51632 48872
rect 51626 48832 51632 48844
rect 51684 48832 51690 48884
rect 47578 48804 47584 48816
rect 45833 48767 45891 48773
rect 45940 48776 47072 48804
rect 47539 48776 47584 48804
rect 43901 48739 43959 48745
rect 43901 48705 43913 48739
rect 43947 48705 43959 48739
rect 43901 48699 43959 48705
rect 43165 48671 43223 48677
rect 43165 48637 43177 48671
rect 43211 48637 43223 48671
rect 43916 48668 43944 48699
rect 45094 48696 45100 48748
rect 45152 48736 45158 48748
rect 45940 48736 45968 48776
rect 46198 48736 46204 48748
rect 45152 48708 45968 48736
rect 46159 48708 46204 48736
rect 45152 48696 45158 48708
rect 46198 48696 46204 48708
rect 46256 48696 46262 48748
rect 47044 48745 47072 48776
rect 47578 48764 47584 48776
rect 47636 48764 47642 48816
rect 47670 48764 47676 48816
rect 47728 48804 47734 48816
rect 50525 48807 50583 48813
rect 50525 48804 50537 48807
rect 47728 48776 50537 48804
rect 47728 48764 47734 48776
rect 48884 48745 48912 48776
rect 50525 48773 50537 48776
rect 50571 48773 50583 48807
rect 50525 48767 50583 48773
rect 46753 48739 46811 48745
rect 46753 48705 46765 48739
rect 46799 48705 46811 48739
rect 46753 48699 46811 48705
rect 47029 48739 47087 48745
rect 47029 48705 47041 48739
rect 47075 48705 47087 48739
rect 47029 48699 47087 48705
rect 48869 48739 48927 48745
rect 48869 48705 48881 48739
rect 48915 48705 48927 48739
rect 48869 48699 48927 48705
rect 49605 48739 49663 48745
rect 49605 48705 49617 48739
rect 49651 48705 49663 48739
rect 49605 48699 49663 48705
rect 46768 48668 46796 48699
rect 47578 48668 47584 48680
rect 43916 48640 45784 48668
rect 46768 48640 47584 48668
rect 43165 48631 43223 48637
rect 40037 48603 40095 48609
rect 40037 48569 40049 48603
rect 40083 48600 40095 48603
rect 41414 48600 41420 48612
rect 40083 48572 41420 48600
rect 40083 48569 40095 48572
rect 40037 48563 40095 48569
rect 41414 48560 41420 48572
rect 41472 48560 41478 48612
rect 45646 48600 45652 48612
rect 45607 48572 45652 48600
rect 45646 48560 45652 48572
rect 45704 48560 45710 48612
rect 45756 48600 45784 48640
rect 47578 48628 47584 48640
rect 47636 48628 47642 48680
rect 49620 48668 49648 48699
rect 50154 48696 50160 48748
rect 50212 48736 50218 48748
rect 50341 48739 50399 48745
rect 50341 48736 50353 48739
rect 50212 48708 50353 48736
rect 50212 48696 50218 48708
rect 50341 48705 50353 48708
rect 50387 48705 50399 48739
rect 50341 48699 50399 48705
rect 51350 48696 51356 48748
rect 51408 48736 51414 48748
rect 51445 48739 51503 48745
rect 51445 48736 51457 48739
rect 51408 48708 51457 48736
rect 51408 48696 51414 48708
rect 51445 48705 51457 48708
rect 51491 48705 51503 48739
rect 51445 48699 51503 48705
rect 51368 48668 51396 48696
rect 49620 48640 51396 48668
rect 45756 48572 47808 48600
rect 40678 48532 40684 48544
rect 39868 48504 40684 48532
rect 38657 48495 38715 48501
rect 40678 48492 40684 48504
rect 40736 48492 40742 48544
rect 40773 48535 40831 48541
rect 40773 48501 40785 48535
rect 40819 48532 40831 48535
rect 40954 48532 40960 48544
rect 40819 48504 40960 48532
rect 40819 48501 40831 48504
rect 40773 48495 40831 48501
rect 40954 48492 40960 48504
rect 41012 48492 41018 48544
rect 45186 48492 45192 48544
rect 45244 48532 45250 48544
rect 46198 48532 46204 48544
rect 45244 48504 46204 48532
rect 45244 48492 45250 48504
rect 46198 48492 46204 48504
rect 46256 48492 46262 48544
rect 46753 48535 46811 48541
rect 46753 48501 46765 48535
rect 46799 48532 46811 48535
rect 47026 48532 47032 48544
rect 46799 48504 47032 48532
rect 46799 48501 46811 48504
rect 46753 48495 46811 48501
rect 47026 48492 47032 48504
rect 47084 48492 47090 48544
rect 47780 48541 47808 48572
rect 47765 48535 47823 48541
rect 47765 48501 47777 48535
rect 47811 48501 47823 48535
rect 47946 48532 47952 48544
rect 47907 48504 47952 48532
rect 47765 48495 47823 48501
rect 47946 48492 47952 48504
rect 48004 48492 48010 48544
rect 48961 48535 49019 48541
rect 48961 48501 48973 48535
rect 49007 48532 49019 48535
rect 49418 48532 49424 48544
rect 49007 48504 49424 48532
rect 49007 48501 49019 48504
rect 48961 48495 49019 48501
rect 49418 48492 49424 48504
rect 49476 48492 49482 48544
rect 49694 48532 49700 48544
rect 49655 48504 49700 48532
rect 49694 48492 49700 48504
rect 49752 48492 49758 48544
rect 1104 48442 68816 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 65654 48442
rect 65706 48390 65718 48442
rect 65770 48390 65782 48442
rect 65834 48390 65846 48442
rect 65898 48390 65910 48442
rect 65962 48390 68816 48442
rect 1104 48368 68816 48390
rect 19794 48328 19800 48340
rect 19755 48300 19800 48328
rect 19794 48288 19800 48300
rect 19852 48288 19858 48340
rect 19978 48328 19984 48340
rect 19939 48300 19984 48328
rect 19978 48288 19984 48300
rect 20036 48288 20042 48340
rect 32692 48300 32996 48328
rect 33704 48314 34100 48328
rect 32692 48272 32720 48300
rect 32968 48272 32996 48300
rect 33545 48300 34100 48314
rect 33545 48286 33732 48300
rect 29362 48260 29368 48272
rect 26206 48232 29368 48260
rect 20438 48192 20444 48204
rect 14476 48164 15700 48192
rect 20399 48164 20444 48192
rect 14476 48136 14504 48164
rect 1670 48084 1676 48136
rect 1728 48124 1734 48136
rect 1949 48127 2007 48133
rect 1949 48124 1961 48127
rect 1728 48096 1961 48124
rect 1728 48084 1734 48096
rect 1949 48093 1961 48096
rect 1995 48093 2007 48127
rect 1949 48087 2007 48093
rect 12897 48127 12955 48133
rect 12897 48093 12909 48127
rect 12943 48124 12955 48127
rect 13354 48124 13360 48136
rect 12943 48096 13360 48124
rect 12943 48093 12955 48096
rect 12897 48087 12955 48093
rect 13354 48084 13360 48096
rect 13412 48084 13418 48136
rect 14458 48124 14464 48136
rect 14371 48096 14464 48124
rect 14458 48084 14464 48096
rect 14516 48084 14522 48136
rect 15197 48127 15255 48133
rect 15197 48093 15209 48127
rect 15243 48124 15255 48127
rect 15286 48124 15292 48136
rect 15243 48096 15292 48124
rect 15243 48093 15255 48096
rect 15197 48087 15255 48093
rect 15286 48084 15292 48096
rect 15344 48084 15350 48136
rect 15672 48133 15700 48164
rect 20438 48152 20444 48164
rect 20496 48152 20502 48204
rect 15657 48127 15715 48133
rect 15657 48093 15669 48127
rect 15703 48093 15715 48127
rect 15657 48087 15715 48093
rect 16485 48127 16543 48133
rect 16485 48093 16497 48127
rect 16531 48124 16543 48127
rect 16758 48124 16764 48136
rect 16531 48096 16764 48124
rect 16531 48093 16543 48096
rect 16485 48087 16543 48093
rect 16758 48084 16764 48096
rect 16816 48084 16822 48136
rect 17221 48127 17279 48133
rect 17221 48093 17233 48127
rect 17267 48124 17279 48127
rect 17402 48124 17408 48136
rect 17267 48096 17408 48124
rect 17267 48093 17279 48096
rect 17221 48087 17279 48093
rect 17402 48084 17408 48096
rect 17460 48084 17466 48136
rect 20714 48133 20720 48136
rect 20708 48124 20720 48133
rect 20675 48096 20720 48124
rect 20708 48087 20720 48096
rect 20714 48084 20720 48087
rect 20772 48084 20778 48136
rect 23201 48127 23259 48133
rect 23201 48093 23213 48127
rect 23247 48093 23259 48127
rect 23201 48087 23259 48093
rect 15749 48059 15807 48065
rect 15749 48025 15761 48059
rect 15795 48056 15807 48059
rect 17954 48056 17960 48068
rect 15795 48028 17960 48056
rect 15795 48025 15807 48028
rect 15749 48019 15807 48025
rect 17954 48016 17960 48028
rect 18012 48016 18018 48068
rect 18046 48016 18052 48068
rect 18104 48056 18110 48068
rect 19613 48059 19671 48065
rect 19613 48056 19625 48059
rect 18104 48028 19625 48056
rect 18104 48016 18110 48028
rect 19613 48025 19625 48028
rect 19659 48056 19671 48059
rect 23216 48056 23244 48087
rect 23290 48084 23296 48136
rect 23348 48124 23354 48136
rect 23348 48096 24256 48124
rect 23348 48084 23354 48096
rect 23658 48056 23664 48068
rect 19659 48028 21864 48056
rect 23216 48028 23664 48056
rect 19659 48025 19671 48028
rect 19613 48019 19671 48025
rect 12710 47988 12716 48000
rect 12671 47960 12716 47988
rect 12710 47948 12716 47960
rect 12768 47948 12774 48000
rect 14182 47948 14188 48000
rect 14240 47988 14246 48000
rect 14461 47991 14519 47997
rect 14461 47988 14473 47991
rect 14240 47960 14473 47988
rect 14240 47948 14246 47960
rect 14461 47957 14473 47960
rect 14507 47957 14519 47991
rect 15010 47988 15016 48000
rect 14971 47960 15016 47988
rect 14461 47951 14519 47957
rect 15010 47948 15016 47960
rect 15068 47948 15074 48000
rect 16298 47948 16304 48000
rect 16356 47988 16362 48000
rect 16485 47991 16543 47997
rect 16485 47988 16497 47991
rect 16356 47960 16497 47988
rect 16356 47948 16362 47960
rect 16485 47957 16497 47960
rect 16531 47957 16543 47991
rect 17034 47988 17040 48000
rect 16995 47960 17040 47988
rect 16485 47951 16543 47957
rect 17034 47948 17040 47960
rect 17092 47948 17098 48000
rect 19823 47991 19881 47997
rect 19823 47957 19835 47991
rect 19869 47988 19881 47991
rect 20162 47988 20168 48000
rect 19869 47960 20168 47988
rect 19869 47957 19881 47960
rect 19823 47951 19881 47957
rect 20162 47948 20168 47960
rect 20220 47948 20226 48000
rect 21836 47997 21864 48028
rect 23658 48016 23664 48028
rect 23716 48016 23722 48068
rect 24228 48056 24256 48096
rect 24302 48084 24308 48136
rect 24360 48124 24366 48136
rect 24397 48127 24455 48133
rect 24397 48124 24409 48127
rect 24360 48096 24409 48124
rect 24360 48084 24366 48096
rect 24397 48093 24409 48096
rect 24443 48093 24455 48127
rect 24397 48087 24455 48093
rect 24664 48127 24722 48133
rect 24664 48093 24676 48127
rect 24710 48124 24722 48127
rect 25406 48124 25412 48136
rect 24710 48096 25412 48124
rect 24710 48093 24722 48096
rect 24664 48087 24722 48093
rect 25406 48084 25412 48096
rect 25464 48084 25470 48136
rect 26206 48124 26234 48232
rect 29362 48220 29368 48232
rect 29420 48260 29426 48272
rect 30282 48260 30288 48272
rect 29420 48232 30288 48260
rect 29420 48220 29426 48232
rect 30282 48220 30288 48232
rect 30340 48220 30346 48272
rect 30374 48220 30380 48272
rect 30432 48260 30438 48272
rect 31570 48260 31576 48272
rect 30432 48232 31576 48260
rect 30432 48220 30438 48232
rect 31570 48220 31576 48232
rect 31628 48260 31634 48272
rect 32217 48263 32275 48269
rect 32217 48260 32229 48263
rect 31628 48232 32229 48260
rect 31628 48220 31634 48232
rect 32217 48229 32229 48232
rect 32263 48229 32275 48263
rect 32217 48223 32275 48229
rect 32674 48220 32680 48272
rect 32732 48220 32738 48272
rect 32858 48260 32864 48272
rect 32819 48232 32864 48260
rect 32858 48220 32864 48232
rect 32916 48220 32922 48272
rect 32950 48220 32956 48272
rect 33008 48220 33014 48272
rect 30392 48192 30420 48220
rect 33545 48192 33573 48286
rect 34072 48260 34100 48300
rect 37200 48300 37504 48328
rect 37200 48260 37228 48300
rect 37366 48260 37372 48272
rect 34072 48232 37228 48260
rect 37327 48232 37372 48260
rect 37366 48220 37372 48232
rect 37424 48220 37430 48272
rect 37476 48260 37504 48300
rect 41322 48288 41328 48340
rect 41380 48328 41386 48340
rect 41601 48331 41659 48337
rect 41601 48328 41613 48331
rect 41380 48300 41613 48328
rect 41380 48288 41386 48300
rect 41601 48297 41613 48300
rect 41647 48328 41659 48331
rect 41874 48328 41880 48340
rect 41647 48300 41880 48328
rect 41647 48297 41659 48300
rect 41601 48291 41659 48297
rect 41874 48288 41880 48300
rect 41932 48288 41938 48340
rect 42720 48300 43668 48328
rect 39482 48260 39488 48272
rect 37476 48232 39488 48260
rect 39482 48220 39488 48232
rect 39540 48220 39546 48272
rect 41782 48260 41788 48272
rect 41743 48232 41788 48260
rect 41782 48220 41788 48232
rect 41840 48220 41846 48272
rect 26344 48164 30420 48192
rect 30484 48164 33573 48192
rect 26344 48133 26372 48164
rect 26068 48096 26234 48124
rect 26329 48127 26387 48133
rect 26068 48056 26096 48096
rect 26329 48093 26341 48127
rect 26375 48093 26387 48127
rect 26329 48087 26387 48093
rect 27341 48127 27399 48133
rect 27341 48093 27353 48127
rect 27387 48124 27399 48127
rect 27522 48124 27528 48136
rect 27387 48096 27528 48124
rect 27387 48093 27399 48096
rect 27341 48087 27399 48093
rect 24228 48028 26096 48056
rect 21821 47991 21879 47997
rect 21821 47957 21833 47991
rect 21867 47957 21879 47991
rect 21821 47951 21879 47957
rect 23290 47948 23296 48000
rect 23348 47988 23354 48000
rect 23477 47991 23535 47997
rect 23477 47988 23489 47991
rect 23348 47960 23489 47988
rect 23348 47948 23354 47960
rect 23477 47957 23489 47960
rect 23523 47957 23535 47991
rect 23477 47951 23535 47957
rect 24854 47948 24860 48000
rect 24912 47988 24918 48000
rect 25777 47991 25835 47997
rect 25777 47988 25789 47991
rect 24912 47960 25789 47988
rect 24912 47948 24918 47960
rect 25777 47957 25789 47960
rect 25823 47957 25835 47991
rect 25777 47951 25835 47957
rect 25866 47948 25872 48000
rect 25924 47988 25930 48000
rect 26344 47988 26372 48087
rect 27522 48084 27528 48096
rect 27580 48084 27586 48136
rect 30484 48133 30512 48164
rect 33686 48152 33692 48204
rect 33744 48192 33750 48204
rect 33873 48195 33931 48201
rect 33744 48164 33789 48192
rect 33744 48152 33750 48164
rect 33873 48161 33885 48195
rect 33919 48161 33931 48195
rect 33873 48155 33931 48161
rect 29733 48127 29791 48133
rect 29733 48093 29745 48127
rect 29779 48124 29791 48127
rect 30469 48127 30527 48133
rect 30469 48124 30481 48127
rect 29779 48096 30481 48124
rect 29779 48093 29791 48096
rect 29733 48087 29791 48093
rect 30469 48093 30481 48096
rect 30515 48093 30527 48127
rect 30469 48087 30527 48093
rect 30558 48084 30564 48136
rect 30616 48124 30622 48136
rect 31297 48127 31355 48133
rect 31297 48124 31309 48127
rect 30616 48096 31309 48124
rect 30616 48084 30622 48096
rect 31297 48093 31309 48096
rect 31343 48093 31355 48127
rect 32674 48124 32680 48136
rect 31297 48087 31355 48093
rect 31404 48096 32680 48124
rect 27430 48016 27436 48068
rect 27488 48056 27494 48068
rect 31404 48056 31432 48096
rect 32674 48084 32680 48096
rect 32732 48084 32738 48136
rect 33134 48124 33140 48136
rect 33095 48096 33140 48124
rect 33134 48084 33140 48096
rect 33192 48084 33198 48136
rect 33597 48127 33655 48133
rect 33597 48124 33609 48127
rect 33520 48096 33609 48124
rect 27488 48028 31432 48056
rect 32033 48059 32091 48065
rect 27488 48016 27494 48028
rect 32033 48025 32045 48059
rect 32079 48056 32091 48059
rect 32490 48056 32496 48068
rect 32079 48028 32496 48056
rect 32079 48025 32091 48028
rect 32033 48019 32091 48025
rect 32490 48016 32496 48028
rect 32548 48016 32554 48068
rect 32861 48059 32919 48065
rect 32861 48025 32873 48059
rect 32907 48056 32919 48059
rect 33226 48056 33232 48068
rect 32907 48028 33232 48056
rect 32907 48025 32919 48028
rect 32861 48019 32919 48025
rect 33226 48016 33232 48028
rect 33284 48016 33290 48068
rect 25924 47960 26372 47988
rect 26421 47991 26479 47997
rect 25924 47948 25930 47960
rect 26421 47957 26433 47991
rect 26467 47988 26479 47991
rect 26510 47988 26516 48000
rect 26467 47960 26516 47988
rect 26467 47957 26479 47960
rect 26421 47951 26479 47957
rect 26510 47948 26516 47960
rect 26568 47948 26574 48000
rect 27154 47988 27160 48000
rect 27115 47960 27160 47988
rect 27154 47948 27160 47960
rect 27212 47948 27218 48000
rect 29178 47948 29184 48000
rect 29236 47988 29242 48000
rect 29825 47991 29883 47997
rect 29825 47988 29837 47991
rect 29236 47960 29837 47988
rect 29236 47948 29242 47960
rect 29825 47957 29837 47960
rect 29871 47957 29883 47991
rect 29825 47951 29883 47957
rect 30190 47948 30196 48000
rect 30248 47988 30254 48000
rect 30561 47991 30619 47997
rect 30561 47988 30573 47991
rect 30248 47960 30573 47988
rect 30248 47948 30254 47960
rect 30561 47957 30573 47960
rect 30607 47957 30619 47991
rect 31110 47988 31116 48000
rect 31071 47960 31116 47988
rect 30561 47951 30619 47957
rect 31110 47948 31116 47960
rect 31168 47948 31174 48000
rect 32950 47948 32956 48000
rect 33008 47988 33014 48000
rect 33045 47991 33103 47997
rect 33045 47988 33057 47991
rect 33008 47960 33057 47988
rect 33008 47948 33014 47960
rect 33045 47957 33057 47960
rect 33091 47988 33103 47991
rect 33520 47988 33548 48096
rect 33597 48093 33609 48096
rect 33643 48093 33655 48127
rect 33888 48124 33916 48155
rect 33962 48152 33968 48204
rect 34020 48192 34026 48204
rect 40126 48192 40132 48204
rect 34020 48164 40132 48192
rect 34020 48152 34026 48164
rect 40126 48152 40132 48164
rect 40184 48152 40190 48204
rect 40313 48195 40371 48201
rect 40313 48161 40325 48195
rect 40359 48192 40371 48195
rect 41506 48192 41512 48204
rect 40359 48164 41512 48192
rect 40359 48161 40371 48164
rect 40313 48155 40371 48161
rect 41506 48152 41512 48164
rect 41564 48192 41570 48204
rect 41690 48192 41696 48204
rect 41564 48164 41696 48192
rect 41564 48152 41570 48164
rect 41690 48152 41696 48164
rect 41748 48192 41754 48204
rect 42720 48192 42748 48300
rect 43073 48263 43131 48269
rect 43073 48229 43085 48263
rect 43119 48260 43131 48263
rect 43162 48260 43168 48272
rect 43119 48232 43168 48260
rect 43119 48229 43131 48232
rect 43073 48223 43131 48229
rect 43162 48220 43168 48232
rect 43220 48220 43226 48272
rect 43640 48260 43668 48300
rect 43714 48288 43720 48340
rect 43772 48328 43778 48340
rect 43809 48331 43867 48337
rect 43809 48328 43821 48331
rect 43772 48300 43821 48328
rect 43772 48288 43778 48300
rect 43809 48297 43821 48300
rect 43855 48297 43867 48331
rect 43809 48291 43867 48297
rect 43898 48288 43904 48340
rect 43956 48328 43962 48340
rect 45373 48331 45431 48337
rect 45373 48328 45385 48331
rect 43956 48300 45385 48328
rect 43956 48288 43962 48300
rect 45373 48297 45385 48300
rect 45419 48297 45431 48331
rect 45373 48291 45431 48297
rect 45833 48331 45891 48337
rect 45833 48297 45845 48331
rect 45879 48328 45891 48331
rect 46014 48328 46020 48340
rect 45879 48300 46020 48328
rect 45879 48297 45891 48300
rect 45833 48291 45891 48297
rect 46014 48288 46020 48300
rect 46072 48288 46078 48340
rect 43916 48260 43944 48288
rect 47026 48260 47032 48272
rect 43640 48232 43944 48260
rect 46987 48232 47032 48260
rect 47026 48220 47032 48232
rect 47084 48220 47090 48272
rect 49237 48263 49295 48269
rect 49237 48229 49249 48263
rect 49283 48260 49295 48263
rect 49283 48232 49648 48260
rect 49283 48229 49295 48232
rect 49237 48223 49295 48229
rect 41748 48164 42748 48192
rect 41748 48152 41754 48164
rect 43254 48152 43260 48204
rect 43312 48192 43318 48204
rect 43533 48195 43591 48201
rect 43533 48192 43545 48195
rect 43312 48164 43545 48192
rect 43312 48152 43318 48164
rect 43533 48161 43545 48164
rect 43579 48161 43591 48195
rect 43533 48155 43591 48161
rect 44361 48195 44419 48201
rect 44361 48161 44373 48195
rect 44407 48192 44419 48195
rect 45002 48192 45008 48204
rect 44407 48164 45008 48192
rect 44407 48161 44419 48164
rect 44361 48155 44419 48161
rect 45002 48152 45008 48164
rect 45060 48152 45066 48204
rect 45557 48195 45615 48201
rect 45557 48192 45569 48195
rect 45112 48164 45569 48192
rect 34422 48124 34428 48136
rect 33888 48096 34428 48124
rect 33597 48087 33655 48093
rect 34422 48084 34428 48096
rect 34480 48084 34486 48136
rect 35618 48084 35624 48136
rect 35676 48124 35682 48136
rect 36170 48124 36176 48136
rect 35676 48096 36176 48124
rect 35676 48084 35682 48096
rect 36170 48084 36176 48096
rect 36228 48084 36234 48136
rect 37093 48127 37151 48133
rect 37093 48093 37105 48127
rect 37139 48093 37151 48127
rect 37093 48087 37151 48093
rect 37185 48127 37243 48133
rect 37185 48093 37197 48127
rect 37231 48124 37243 48127
rect 37274 48124 37280 48136
rect 37231 48096 37280 48124
rect 37231 48093 37243 48096
rect 37185 48087 37243 48093
rect 33870 48056 33876 48068
rect 33831 48028 33876 48056
rect 33870 48016 33876 48028
rect 33928 48016 33934 48068
rect 37108 48056 37136 48087
rect 37274 48084 37280 48096
rect 37332 48084 37338 48136
rect 40034 48124 40040 48136
rect 39995 48096 40040 48124
rect 40034 48084 40040 48096
rect 40092 48084 40098 48136
rect 40218 48124 40224 48136
rect 40179 48096 40224 48124
rect 40218 48084 40224 48096
rect 40276 48084 40282 48136
rect 44266 48124 44272 48136
rect 40328 48096 43576 48124
rect 44227 48096 44272 48124
rect 37918 48056 37924 48068
rect 37108 48028 37924 48056
rect 37918 48016 37924 48028
rect 37976 48016 37982 48068
rect 38010 48016 38016 48068
rect 38068 48056 38074 48068
rect 40328 48056 40356 48096
rect 38068 48028 40356 48056
rect 38068 48016 38074 48028
rect 40678 48016 40684 48068
rect 40736 48056 40742 48068
rect 41322 48056 41328 48068
rect 40736 48028 41328 48056
rect 40736 48016 40742 48028
rect 41322 48016 41328 48028
rect 41380 48056 41386 48068
rect 41417 48059 41475 48065
rect 41417 48056 41429 48059
rect 41380 48028 41429 48056
rect 41380 48016 41386 48028
rect 41417 48025 41429 48028
rect 41463 48025 41475 48059
rect 41417 48019 41475 48025
rect 41598 48016 41604 48068
rect 41656 48065 41662 48068
rect 41656 48059 41675 48065
rect 41663 48025 41675 48059
rect 43070 48056 43076 48068
rect 43031 48028 43076 48056
rect 41656 48019 41675 48025
rect 41656 48016 41662 48019
rect 43070 48016 43076 48028
rect 43128 48016 43134 48068
rect 43548 48056 43576 48096
rect 44266 48084 44272 48096
rect 44324 48084 44330 48136
rect 44450 48124 44456 48136
rect 44411 48096 44456 48124
rect 44450 48084 44456 48096
rect 44508 48084 44514 48136
rect 44910 48084 44916 48136
rect 44968 48124 44974 48136
rect 45112 48124 45140 48164
rect 45557 48161 45569 48164
rect 45603 48161 45615 48195
rect 45557 48155 45615 48161
rect 47118 48152 47124 48204
rect 47176 48192 47182 48204
rect 47213 48195 47271 48201
rect 47213 48192 47225 48195
rect 47176 48164 47225 48192
rect 47176 48152 47182 48164
rect 47213 48161 47225 48164
rect 47259 48161 47271 48195
rect 47213 48155 47271 48161
rect 48516 48164 49280 48192
rect 45278 48124 45284 48136
rect 44968 48096 45140 48124
rect 45239 48096 45284 48124
rect 44968 48084 44974 48096
rect 45278 48084 45284 48096
rect 45336 48084 45342 48136
rect 45462 48084 45468 48136
rect 45520 48124 45526 48136
rect 46937 48127 46995 48133
rect 45520 48096 46888 48124
rect 45520 48084 45526 48096
rect 45646 48056 45652 48068
rect 43548 48028 45652 48056
rect 45646 48016 45652 48028
rect 45704 48016 45710 48068
rect 46860 48056 46888 48096
rect 46937 48093 46949 48127
rect 46983 48124 46995 48127
rect 47946 48124 47952 48136
rect 46983 48096 47952 48124
rect 46983 48093 46995 48096
rect 46937 48087 46995 48093
rect 47946 48084 47952 48096
rect 48004 48084 48010 48136
rect 48516 48133 48544 48164
rect 48501 48127 48559 48133
rect 48501 48124 48513 48127
rect 48056 48096 48513 48124
rect 48056 48056 48084 48096
rect 48501 48093 48513 48096
rect 48547 48093 48559 48127
rect 48501 48087 48559 48093
rect 48682 48084 48688 48136
rect 48740 48124 48746 48136
rect 48777 48127 48835 48133
rect 48777 48124 48789 48127
rect 48740 48096 48789 48124
rect 48740 48084 48746 48096
rect 48777 48093 48789 48096
rect 48823 48093 48835 48127
rect 48777 48087 48835 48093
rect 46860 48028 48084 48056
rect 48317 48059 48375 48065
rect 48317 48025 48329 48059
rect 48363 48056 48375 48059
rect 49142 48056 49148 48068
rect 48363 48028 49148 48056
rect 48363 48025 48375 48028
rect 48317 48019 48375 48025
rect 49142 48016 49148 48028
rect 49200 48016 49206 48068
rect 49252 48065 49280 48164
rect 49418 48124 49424 48136
rect 49379 48096 49424 48124
rect 49418 48084 49424 48096
rect 49476 48084 49482 48136
rect 49513 48127 49571 48133
rect 49513 48093 49525 48127
rect 49559 48093 49571 48127
rect 49620 48124 49648 48232
rect 49694 48152 49700 48204
rect 49752 48192 49758 48204
rect 50157 48195 50215 48201
rect 50157 48192 50169 48195
rect 49752 48164 50169 48192
rect 49752 48152 49758 48164
rect 50157 48161 50169 48164
rect 50203 48161 50215 48195
rect 50157 48155 50215 48161
rect 50413 48127 50471 48133
rect 50413 48124 50425 48127
rect 49620 48096 50425 48124
rect 49513 48087 49571 48093
rect 50413 48093 50425 48096
rect 50459 48093 50471 48127
rect 50413 48087 50471 48093
rect 49237 48059 49295 48065
rect 49237 48025 49249 48059
rect 49283 48025 49295 48059
rect 49528 48056 49556 48087
rect 67726 48056 67732 48068
rect 49237 48019 49295 48025
rect 49344 48028 49556 48056
rect 67687 48028 67732 48056
rect 39850 47988 39856 48000
rect 33091 47960 33548 47988
rect 39811 47960 39856 47988
rect 33091 47957 33103 47960
rect 33045 47951 33103 47957
rect 39850 47948 39856 47960
rect 39908 47948 39914 48000
rect 42610 47948 42616 48000
rect 42668 47988 42674 48000
rect 43625 47991 43683 47997
rect 43625 47988 43637 47991
rect 42668 47960 43637 47988
rect 42668 47948 42674 47960
rect 43625 47957 43637 47960
rect 43671 47957 43683 47991
rect 47210 47988 47216 48000
rect 47171 47960 47216 47988
rect 43625 47951 43683 47957
rect 47210 47948 47216 47960
rect 47268 47948 47274 48000
rect 47486 47948 47492 48000
rect 47544 47988 47550 48000
rect 48685 47991 48743 47997
rect 48685 47988 48697 47991
rect 47544 47960 48697 47988
rect 47544 47948 47550 47960
rect 48685 47957 48697 47960
rect 48731 47988 48743 47991
rect 49344 47988 49372 48028
rect 67726 48016 67732 48028
rect 67784 48016 67790 48068
rect 48731 47960 49372 47988
rect 48731 47957 48743 47960
rect 48685 47951 48743 47957
rect 50154 47948 50160 48000
rect 50212 47988 50218 48000
rect 51537 47991 51595 47997
rect 51537 47988 51549 47991
rect 50212 47960 51549 47988
rect 50212 47948 50218 47960
rect 51537 47957 51549 47960
rect 51583 47957 51595 47991
rect 67818 47988 67824 48000
rect 67779 47960 67824 47988
rect 51537 47951 51595 47957
rect 67818 47948 67824 47960
rect 67876 47948 67882 48000
rect 1104 47898 68816 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 68816 47898
rect 1104 47824 68816 47846
rect 17402 47784 17408 47796
rect 17363 47756 17408 47784
rect 17402 47744 17408 47756
rect 17460 47744 17466 47796
rect 17954 47744 17960 47796
rect 18012 47784 18018 47796
rect 24302 47784 24308 47796
rect 18012 47756 22324 47784
rect 24263 47756 24308 47784
rect 18012 47744 18018 47756
rect 12428 47719 12486 47725
rect 12428 47685 12440 47719
rect 12474 47716 12486 47719
rect 12710 47716 12716 47728
rect 12474 47688 12716 47716
rect 12474 47685 12486 47688
rect 12428 47679 12486 47685
rect 12710 47676 12716 47688
rect 12768 47676 12774 47728
rect 14452 47719 14510 47725
rect 14452 47685 14464 47719
rect 14498 47716 14510 47719
rect 15010 47716 15016 47728
rect 14498 47688 15016 47716
rect 14498 47685 14510 47688
rect 14452 47679 14510 47685
rect 15010 47676 15016 47688
rect 15068 47676 15074 47728
rect 1670 47648 1676 47660
rect 1631 47620 1676 47648
rect 1670 47608 1676 47620
rect 1728 47608 1734 47660
rect 14182 47648 14188 47660
rect 14143 47620 14188 47648
rect 14182 47608 14188 47620
rect 14240 47608 14246 47660
rect 17221 47651 17279 47657
rect 17221 47617 17233 47651
rect 17267 47648 17279 47651
rect 17310 47648 17316 47660
rect 17267 47620 17316 47648
rect 17267 47617 17279 47620
rect 17221 47611 17279 47617
rect 17310 47608 17316 47620
rect 17368 47608 17374 47660
rect 18046 47648 18052 47660
rect 18007 47620 18052 47648
rect 18046 47608 18052 47620
rect 18104 47608 18110 47660
rect 22296 47657 22324 47756
rect 24302 47744 24308 47756
rect 24360 47744 24366 47796
rect 27522 47784 27528 47796
rect 27483 47756 27528 47784
rect 27522 47744 27528 47756
rect 27580 47744 27586 47796
rect 33778 47784 33784 47796
rect 28276 47756 33784 47784
rect 25866 47716 25872 47728
rect 22388 47688 25872 47716
rect 22281 47651 22339 47657
rect 22281 47617 22293 47651
rect 22327 47617 22339 47651
rect 22281 47611 22339 47617
rect 1857 47583 1915 47589
rect 1857 47549 1869 47583
rect 1903 47580 1915 47583
rect 2406 47580 2412 47592
rect 1903 47552 2412 47580
rect 1903 47549 1915 47552
rect 1857 47543 1915 47549
rect 2406 47540 2412 47552
rect 2464 47540 2470 47592
rect 2774 47580 2780 47592
rect 2735 47552 2780 47580
rect 2774 47540 2780 47552
rect 2832 47540 2838 47592
rect 12158 47580 12164 47592
rect 12119 47552 12164 47580
rect 12158 47540 12164 47552
rect 12216 47540 12222 47592
rect 17037 47583 17095 47589
rect 17037 47549 17049 47583
rect 17083 47580 17095 47583
rect 17678 47580 17684 47592
rect 17083 47552 17684 47580
rect 17083 47549 17095 47552
rect 17037 47543 17095 47549
rect 17678 47540 17684 47552
rect 17736 47580 17742 47592
rect 17865 47583 17923 47589
rect 17865 47580 17877 47583
rect 17736 47552 17877 47580
rect 17736 47540 17742 47552
rect 17865 47549 17877 47552
rect 17911 47549 17923 47583
rect 18785 47583 18843 47589
rect 18785 47580 18797 47583
rect 17865 47543 17923 47549
rect 18156 47552 18797 47580
rect 15562 47512 15568 47524
rect 15475 47484 15568 47512
rect 15562 47472 15568 47484
rect 15620 47512 15626 47524
rect 18156 47512 18184 47552
rect 18785 47549 18797 47552
rect 18831 47549 18843 47583
rect 18785 47543 18843 47549
rect 18874 47540 18880 47592
rect 18932 47589 18938 47592
rect 18932 47583 18960 47589
rect 18948 47549 18960 47583
rect 18932 47543 18960 47549
rect 18932 47540 18938 47543
rect 19058 47540 19064 47592
rect 19116 47580 19122 47592
rect 19116 47552 19161 47580
rect 19116 47540 19122 47552
rect 20990 47540 20996 47592
rect 21048 47580 21054 47592
rect 22388 47580 22416 47688
rect 25866 47676 25872 47688
rect 25924 47676 25930 47728
rect 27798 47716 27804 47728
rect 27264 47688 27804 47716
rect 22548 47651 22606 47657
rect 22548 47617 22560 47651
rect 22594 47648 22606 47651
rect 23106 47648 23112 47660
rect 22594 47620 23112 47648
rect 22594 47617 22606 47620
rect 22548 47611 22606 47617
rect 23106 47608 23112 47620
rect 23164 47608 23170 47660
rect 24302 47648 24308 47660
rect 24263 47620 24308 47648
rect 24302 47608 24308 47620
rect 24360 47608 24366 47660
rect 26234 47608 26240 47660
rect 26292 47648 26298 47660
rect 27264 47657 27292 47688
rect 27798 47676 27804 47688
rect 27856 47716 27862 47728
rect 28169 47719 28227 47725
rect 28169 47716 28181 47719
rect 27856 47688 28181 47716
rect 27856 47676 27862 47688
rect 28169 47685 28181 47688
rect 28215 47685 28227 47719
rect 28169 47679 28227 47685
rect 27249 47651 27307 47657
rect 26292 47620 26337 47648
rect 26292 47608 26298 47620
rect 27249 47617 27261 47651
rect 27295 47617 27307 47651
rect 27249 47611 27307 47617
rect 27341 47651 27399 47657
rect 27341 47617 27353 47651
rect 27387 47648 27399 47651
rect 27430 47648 27436 47660
rect 27387 47620 27436 47648
rect 27387 47617 27399 47620
rect 27341 47611 27399 47617
rect 27430 47608 27436 47620
rect 27488 47608 27494 47660
rect 28276 47648 28304 47756
rect 33778 47744 33784 47756
rect 33836 47744 33842 47796
rect 33962 47744 33968 47796
rect 34020 47784 34026 47796
rect 34977 47787 35035 47793
rect 34977 47784 34989 47787
rect 34020 47756 34989 47784
rect 34020 47744 34026 47756
rect 34977 47753 34989 47756
rect 35023 47753 35035 47787
rect 34977 47747 35035 47753
rect 35434 47744 35440 47796
rect 35492 47784 35498 47796
rect 35802 47784 35808 47796
rect 35492 47756 35808 47784
rect 35492 47744 35498 47756
rect 35802 47744 35808 47756
rect 35860 47744 35866 47796
rect 35986 47744 35992 47796
rect 36044 47784 36050 47796
rect 67818 47784 67824 47796
rect 36044 47756 67824 47784
rect 36044 47744 36050 47756
rect 67818 47744 67824 47756
rect 67876 47744 67882 47796
rect 28534 47716 28540 47728
rect 28495 47688 28540 47716
rect 28534 47676 28540 47688
rect 28592 47676 28598 47728
rect 28905 47719 28963 47725
rect 28905 47685 28917 47719
rect 28951 47716 28963 47719
rect 29086 47716 29092 47728
rect 28951 47688 29092 47716
rect 28951 47685 28963 47688
rect 28905 47679 28963 47685
rect 29086 47676 29092 47688
rect 29144 47676 29150 47728
rect 29273 47719 29331 47725
rect 29273 47685 29285 47719
rect 29319 47685 29331 47719
rect 29273 47679 29331 47685
rect 30460 47719 30518 47725
rect 30460 47685 30472 47719
rect 30506 47716 30518 47719
rect 31110 47716 31116 47728
rect 30506 47688 31116 47716
rect 30506 47685 30518 47688
rect 30460 47679 30518 47685
rect 28442 47648 28448 47660
rect 27908 47620 28304 47648
rect 28403 47620 28448 47648
rect 21048 47552 22416 47580
rect 21048 47540 21054 47552
rect 25866 47540 25872 47592
rect 25924 47580 25930 47592
rect 27908 47580 27936 47620
rect 28442 47608 28448 47620
rect 28500 47608 28506 47660
rect 25924 47552 27936 47580
rect 25924 47540 25930 47552
rect 28902 47540 28908 47592
rect 28960 47540 28966 47592
rect 29288 47580 29316 47679
rect 31110 47676 31116 47688
rect 31168 47676 31174 47728
rect 34698 47716 34704 47728
rect 32600 47688 34704 47716
rect 30190 47648 30196 47660
rect 30151 47620 30196 47648
rect 30190 47608 30196 47620
rect 30248 47608 30254 47660
rect 32600 47657 32628 47688
rect 34698 47676 34704 47688
rect 34756 47676 34762 47728
rect 35526 47716 35532 47728
rect 35084 47688 35532 47716
rect 32858 47657 32864 47660
rect 32585 47651 32643 47657
rect 32585 47617 32597 47651
rect 32631 47617 32643 47651
rect 32852 47648 32864 47657
rect 32819 47620 32864 47648
rect 32585 47611 32643 47617
rect 32852 47611 32864 47620
rect 32858 47608 32864 47611
rect 32916 47608 32922 47660
rect 33134 47608 33140 47660
rect 33192 47648 33198 47660
rect 33192 47620 33640 47648
rect 33192 47608 33198 47620
rect 33612 47580 33640 47620
rect 33778 47608 33784 47660
rect 33836 47648 33842 47660
rect 35084 47657 35112 47688
rect 35526 47676 35532 47688
rect 35584 47716 35590 47728
rect 36081 47719 36139 47725
rect 36081 47716 36093 47719
rect 35584 47688 36093 47716
rect 35584 47676 35590 47688
rect 36081 47685 36093 47688
rect 36127 47685 36139 47719
rect 36081 47679 36139 47685
rect 36354 47676 36360 47728
rect 36412 47716 36418 47728
rect 40865 47719 40923 47725
rect 40865 47716 40877 47719
rect 36412 47688 39160 47716
rect 36412 47676 36418 47688
rect 34793 47651 34851 47657
rect 34793 47648 34805 47651
rect 33836 47620 34805 47648
rect 33836 47608 33842 47620
rect 34793 47617 34805 47620
rect 34839 47617 34851 47651
rect 34793 47611 34851 47617
rect 35069 47651 35127 47657
rect 35069 47617 35081 47651
rect 35115 47617 35127 47651
rect 35069 47611 35127 47617
rect 35618 47608 35624 47660
rect 35676 47648 35682 47660
rect 35713 47651 35771 47657
rect 35713 47648 35725 47651
rect 35676 47620 35725 47648
rect 35676 47608 35682 47620
rect 35713 47617 35725 47620
rect 35759 47617 35771 47651
rect 35713 47611 35771 47617
rect 35897 47651 35955 47657
rect 35897 47617 35909 47651
rect 35943 47617 35955 47651
rect 37826 47648 37832 47660
rect 37787 47620 37832 47648
rect 35897 47611 35955 47617
rect 33686 47580 33692 47592
rect 29288 47552 30236 47580
rect 33612 47552 33692 47580
rect 15620 47484 18184 47512
rect 15620 47472 15626 47484
rect 18230 47472 18236 47524
rect 18288 47512 18294 47524
rect 18509 47515 18567 47521
rect 18509 47512 18521 47515
rect 18288 47484 18521 47512
rect 18288 47472 18294 47484
rect 18509 47481 18521 47484
rect 18555 47481 18567 47515
rect 18509 47475 18567 47481
rect 30208 47456 30236 47552
rect 33686 47540 33692 47552
rect 33744 47580 33750 47592
rect 34330 47580 34336 47592
rect 33744 47552 34336 47580
rect 33744 47540 33750 47552
rect 34330 47540 34336 47552
rect 34388 47540 34394 47592
rect 35529 47515 35587 47521
rect 35529 47481 35541 47515
rect 35575 47512 35587 47515
rect 35618 47512 35624 47524
rect 35575 47484 35624 47512
rect 35575 47481 35587 47484
rect 35529 47475 35587 47481
rect 35618 47472 35624 47484
rect 35676 47472 35682 47524
rect 13538 47444 13544 47456
rect 13451 47416 13544 47444
rect 13538 47404 13544 47416
rect 13596 47444 13602 47456
rect 18874 47444 18880 47456
rect 13596 47416 18880 47444
rect 13596 47404 13602 47416
rect 18874 47404 18880 47416
rect 18932 47404 18938 47456
rect 19705 47447 19763 47453
rect 19705 47413 19717 47447
rect 19751 47444 19763 47447
rect 21082 47444 21088 47456
rect 19751 47416 21088 47444
rect 19751 47413 19763 47416
rect 19705 47407 19763 47413
rect 21082 47404 21088 47416
rect 21140 47404 21146 47456
rect 23658 47444 23664 47456
rect 23571 47416 23664 47444
rect 23658 47404 23664 47416
rect 23716 47444 23722 47456
rect 24762 47444 24768 47456
rect 23716 47416 24768 47444
rect 23716 47404 23722 47416
rect 24762 47404 24768 47416
rect 24820 47404 24826 47456
rect 26329 47447 26387 47453
rect 26329 47413 26341 47447
rect 26375 47444 26387 47447
rect 26418 47444 26424 47456
rect 26375 47416 26424 47444
rect 26375 47413 26387 47416
rect 26329 47407 26387 47413
rect 26418 47404 26424 47416
rect 26476 47404 26482 47456
rect 29454 47444 29460 47456
rect 29415 47416 29460 47444
rect 29454 47404 29460 47416
rect 29512 47404 29518 47456
rect 30190 47404 30196 47456
rect 30248 47444 30254 47456
rect 31573 47447 31631 47453
rect 31573 47444 31585 47447
rect 30248 47416 31585 47444
rect 30248 47404 30254 47416
rect 31573 47413 31585 47416
rect 31619 47413 31631 47447
rect 31573 47407 31631 47413
rect 33594 47404 33600 47456
rect 33652 47444 33658 47456
rect 33965 47447 34023 47453
rect 33965 47444 33977 47447
rect 33652 47416 33977 47444
rect 33652 47404 33658 47416
rect 33965 47413 33977 47416
rect 34011 47413 34023 47447
rect 34606 47444 34612 47456
rect 34567 47416 34612 47444
rect 33965 47407 34023 47413
rect 34606 47404 34612 47416
rect 34664 47404 34670 47456
rect 34790 47404 34796 47456
rect 34848 47444 34854 47456
rect 35434 47444 35440 47456
rect 34848 47416 35440 47444
rect 34848 47404 34854 47416
rect 35434 47404 35440 47416
rect 35492 47444 35498 47456
rect 35912 47444 35940 47611
rect 37826 47608 37832 47620
rect 37884 47608 37890 47660
rect 39025 47651 39083 47657
rect 39025 47617 39037 47651
rect 39071 47617 39083 47651
rect 39025 47611 39083 47617
rect 35492 47416 35940 47444
rect 38013 47447 38071 47453
rect 35492 47404 35498 47416
rect 38013 47413 38025 47447
rect 38059 47444 38071 47447
rect 38746 47444 38752 47456
rect 38059 47416 38752 47444
rect 38059 47413 38071 47416
rect 38013 47407 38071 47413
rect 38746 47404 38752 47416
rect 38804 47404 38810 47456
rect 39040 47444 39068 47611
rect 39132 47512 39160 47688
rect 39408 47688 40877 47716
rect 39408 47660 39436 47688
rect 40865 47685 40877 47688
rect 40911 47685 40923 47719
rect 42610 47716 42616 47728
rect 40865 47679 40923 47685
rect 41064 47688 42616 47716
rect 39390 47648 39396 47660
rect 39351 47620 39396 47648
rect 39390 47608 39396 47620
rect 39448 47608 39454 47660
rect 39761 47651 39819 47657
rect 39761 47617 39773 47651
rect 39807 47648 39819 47651
rect 39942 47648 39948 47660
rect 39807 47620 39948 47648
rect 39807 47617 39819 47620
rect 39761 47611 39819 47617
rect 39942 47608 39948 47620
rect 40000 47648 40006 47660
rect 40681 47651 40739 47657
rect 40681 47648 40693 47651
rect 40000 47620 40693 47648
rect 40000 47608 40006 47620
rect 40681 47617 40693 47620
rect 40727 47617 40739 47651
rect 40954 47648 40960 47660
rect 40915 47620 40960 47648
rect 40681 47611 40739 47617
rect 39666 47540 39672 47592
rect 39724 47580 39730 47592
rect 39853 47583 39911 47589
rect 39853 47580 39865 47583
rect 39724 47552 39865 47580
rect 39724 47540 39730 47552
rect 39853 47549 39865 47552
rect 39899 47549 39911 47583
rect 40696 47580 40724 47611
rect 40954 47608 40960 47620
rect 41012 47608 41018 47660
rect 41064 47580 41092 47688
rect 42610 47676 42616 47688
rect 42668 47676 42674 47728
rect 43254 47716 43260 47728
rect 43215 47688 43260 47716
rect 43254 47676 43260 47688
rect 43312 47676 43318 47728
rect 47946 47676 47952 47728
rect 48004 47716 48010 47728
rect 48317 47719 48375 47725
rect 48317 47716 48329 47719
rect 48004 47688 48329 47716
rect 48004 47676 48010 47688
rect 48317 47685 48329 47688
rect 48363 47685 48375 47719
rect 48682 47716 48688 47728
rect 48643 47688 48688 47716
rect 48317 47679 48375 47685
rect 48682 47676 48688 47688
rect 48740 47676 48746 47728
rect 49142 47676 49148 47728
rect 49200 47716 49206 47728
rect 49694 47716 49700 47728
rect 49200 47688 49700 47716
rect 49200 47676 49206 47688
rect 49694 47676 49700 47688
rect 49752 47676 49758 47728
rect 50154 47676 50160 47728
rect 50212 47716 50218 47728
rect 50212 47688 50476 47716
rect 50212 47676 50218 47688
rect 41414 47608 41420 47660
rect 41472 47648 41478 47660
rect 41601 47651 41659 47657
rect 41472 47620 41517 47648
rect 41472 47608 41478 47620
rect 41601 47617 41613 47651
rect 41647 47617 41659 47651
rect 42628 47648 42656 47676
rect 43717 47651 43775 47657
rect 43717 47648 43729 47651
rect 42628 47620 43729 47648
rect 41601 47611 41659 47617
rect 43717 47617 43729 47620
rect 43763 47617 43775 47651
rect 44910 47648 44916 47660
rect 43717 47611 43775 47617
rect 43916 47620 44916 47648
rect 41616 47580 41644 47611
rect 40696 47552 41092 47580
rect 41156 47552 41644 47580
rect 39853 47543 39911 47549
rect 40129 47515 40187 47521
rect 40129 47512 40141 47515
rect 39132 47484 40141 47512
rect 40129 47481 40141 47484
rect 40175 47481 40187 47515
rect 40129 47475 40187 47481
rect 40954 47472 40960 47524
rect 41012 47512 41018 47524
rect 41156 47512 41184 47552
rect 43070 47540 43076 47592
rect 43128 47580 43134 47592
rect 43622 47580 43628 47592
rect 43128 47552 43628 47580
rect 43128 47540 43134 47552
rect 43622 47540 43628 47552
rect 43680 47540 43686 47592
rect 41012 47484 41184 47512
rect 41012 47472 41018 47484
rect 41322 47472 41328 47524
rect 41380 47512 41386 47524
rect 43916 47521 43944 47620
rect 44910 47608 44916 47620
rect 44968 47608 44974 47660
rect 45189 47651 45247 47657
rect 45189 47617 45201 47651
rect 45235 47648 45247 47651
rect 45646 47648 45652 47660
rect 45235 47620 45652 47648
rect 45235 47617 45247 47620
rect 45189 47611 45247 47617
rect 45646 47608 45652 47620
rect 45704 47608 45710 47660
rect 48501 47651 48559 47657
rect 48501 47617 48513 47651
rect 48547 47648 48559 47651
rect 48590 47648 48596 47660
rect 48547 47620 48596 47648
rect 48547 47617 48559 47620
rect 48501 47611 48559 47617
rect 48590 47608 48596 47620
rect 48648 47648 48654 47660
rect 50448 47657 50476 47688
rect 50341 47651 50399 47657
rect 50341 47648 50353 47651
rect 48648 47620 50353 47648
rect 48648 47608 48654 47620
rect 50341 47617 50353 47620
rect 50387 47617 50399 47651
rect 50341 47611 50399 47617
rect 50433 47651 50491 47657
rect 50433 47617 50445 47651
rect 50479 47617 50491 47651
rect 50614 47648 50620 47660
rect 50575 47620 50620 47648
rect 50433 47611 50491 47617
rect 44266 47540 44272 47592
rect 44324 47580 44330 47592
rect 45097 47583 45155 47589
rect 45097 47580 45109 47583
rect 44324 47552 45109 47580
rect 44324 47540 44330 47552
rect 45097 47549 45109 47552
rect 45143 47580 45155 47583
rect 46290 47580 46296 47592
rect 45143 47552 46296 47580
rect 45143 47549 45155 47552
rect 45097 47543 45155 47549
rect 46290 47540 46296 47552
rect 46348 47540 46354 47592
rect 49786 47540 49792 47592
rect 49844 47580 49850 47592
rect 50157 47583 50215 47589
rect 50157 47580 50169 47583
rect 49844 47552 50169 47580
rect 49844 47540 49850 47552
rect 50157 47549 50169 47552
rect 50203 47549 50215 47583
rect 50356 47580 50384 47611
rect 50614 47608 50620 47620
rect 50672 47608 50678 47660
rect 50709 47651 50767 47657
rect 50709 47617 50721 47651
rect 50755 47648 50767 47651
rect 51442 47648 51448 47660
rect 50755 47620 51448 47648
rect 50755 47617 50767 47620
rect 50709 47611 50767 47617
rect 51442 47608 51448 47620
rect 51500 47608 51506 47660
rect 51626 47648 51632 47660
rect 51587 47620 51632 47648
rect 51626 47608 51632 47620
rect 51684 47608 51690 47660
rect 50798 47580 50804 47592
rect 50356 47552 50804 47580
rect 50157 47543 50215 47549
rect 50798 47540 50804 47552
rect 50856 47540 50862 47592
rect 43901 47515 43959 47521
rect 41380 47484 43852 47512
rect 41380 47472 41386 47484
rect 40034 47444 40040 47456
rect 39040 47416 40040 47444
rect 40034 47404 40040 47416
rect 40092 47404 40098 47456
rect 40678 47444 40684 47456
rect 40639 47416 40684 47444
rect 40678 47404 40684 47416
rect 40736 47404 40742 47456
rect 41417 47447 41475 47453
rect 41417 47413 41429 47447
rect 41463 47444 41475 47447
rect 41782 47444 41788 47456
rect 41463 47416 41788 47444
rect 41463 47413 41475 47416
rect 41417 47407 41475 47413
rect 41782 47404 41788 47416
rect 41840 47404 41846 47456
rect 43162 47404 43168 47456
rect 43220 47444 43226 47456
rect 43349 47447 43407 47453
rect 43349 47444 43361 47447
rect 43220 47416 43361 47444
rect 43220 47404 43226 47416
rect 43349 47413 43361 47416
rect 43395 47413 43407 47447
rect 43824 47444 43852 47484
rect 43901 47481 43913 47515
rect 43947 47481 43959 47515
rect 43901 47475 43959 47481
rect 44634 47472 44640 47524
rect 44692 47512 44698 47524
rect 45373 47515 45431 47521
rect 45373 47512 45385 47515
rect 44692 47484 45385 47512
rect 44692 47472 44698 47484
rect 45373 47481 45385 47484
rect 45419 47481 45431 47515
rect 45373 47475 45431 47481
rect 44358 47444 44364 47456
rect 43824 47416 44364 47444
rect 43349 47407 43407 47413
rect 44358 47404 44364 47416
rect 44416 47404 44422 47456
rect 45186 47444 45192 47456
rect 45147 47416 45192 47444
rect 45186 47404 45192 47416
rect 45244 47404 45250 47456
rect 51445 47447 51503 47453
rect 51445 47413 51457 47447
rect 51491 47444 51503 47447
rect 51718 47444 51724 47456
rect 51491 47416 51724 47444
rect 51491 47413 51503 47416
rect 51445 47407 51503 47413
rect 51718 47404 51724 47416
rect 51776 47404 51782 47456
rect 1104 47354 68816 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 65654 47354
rect 65706 47302 65718 47354
rect 65770 47302 65782 47354
rect 65834 47302 65846 47354
rect 65898 47302 65910 47354
rect 65962 47302 68816 47354
rect 1104 47280 68816 47302
rect 2406 47240 2412 47252
rect 2367 47212 2412 47240
rect 2406 47200 2412 47212
rect 2464 47200 2470 47252
rect 12158 47200 12164 47252
rect 12216 47240 12222 47252
rect 12253 47243 12311 47249
rect 12253 47240 12265 47243
rect 12216 47212 12265 47240
rect 12216 47200 12222 47212
rect 12253 47209 12265 47212
rect 12299 47209 12311 47243
rect 13354 47240 13360 47252
rect 13315 47212 13360 47240
rect 12253 47203 12311 47209
rect 13354 47200 13360 47212
rect 13412 47200 13418 47252
rect 15286 47240 15292 47252
rect 15247 47212 15292 47240
rect 15286 47200 15292 47212
rect 15344 47200 15350 47252
rect 17678 47240 17684 47252
rect 17639 47212 17684 47240
rect 17678 47200 17684 47212
rect 17736 47200 17742 47252
rect 23106 47240 23112 47252
rect 23067 47212 23112 47240
rect 23106 47200 23112 47212
rect 23164 47200 23170 47252
rect 27798 47240 27804 47252
rect 27759 47212 27804 47240
rect 27798 47200 27804 47212
rect 27856 47200 27862 47252
rect 30374 47240 30380 47252
rect 30335 47212 30380 47240
rect 30374 47200 30380 47212
rect 30432 47200 30438 47252
rect 30558 47240 30564 47252
rect 30519 47212 30564 47240
rect 30558 47200 30564 47212
rect 30616 47200 30622 47252
rect 32950 47200 32956 47252
rect 33008 47240 33014 47252
rect 33962 47240 33968 47252
rect 33008 47212 33968 47240
rect 33008 47200 33014 47212
rect 33962 47200 33968 47212
rect 34020 47200 34026 47252
rect 38010 47240 38016 47252
rect 34072 47212 38016 47240
rect 14090 47172 14096 47184
rect 12636 47144 14096 47172
rect 12636 47048 12664 47144
rect 14090 47132 14096 47144
rect 14148 47132 14154 47184
rect 29917 47175 29975 47181
rect 29917 47141 29929 47175
rect 29963 47172 29975 47175
rect 30282 47172 30288 47184
rect 29963 47144 30288 47172
rect 29963 47141 29975 47144
rect 29917 47135 29975 47141
rect 30282 47132 30288 47144
rect 30340 47172 30346 47184
rect 34072 47172 34100 47212
rect 38010 47200 38016 47212
rect 38068 47200 38074 47252
rect 39390 47200 39396 47252
rect 39448 47240 39454 47252
rect 40037 47243 40095 47249
rect 40037 47240 40049 47243
rect 39448 47212 40049 47240
rect 39448 47200 39454 47212
rect 40037 47209 40049 47212
rect 40083 47209 40095 47243
rect 40218 47240 40224 47252
rect 40179 47212 40224 47240
rect 40037 47203 40095 47209
rect 30340 47144 34100 47172
rect 34149 47175 34207 47181
rect 30340 47132 30346 47144
rect 34149 47141 34161 47175
rect 34195 47172 34207 47175
rect 34790 47172 34796 47184
rect 34195 47144 34796 47172
rect 34195 47141 34207 47144
rect 34149 47135 34207 47141
rect 34790 47132 34796 47144
rect 34848 47132 34854 47184
rect 34977 47175 35035 47181
rect 34977 47141 34989 47175
rect 35023 47172 35035 47175
rect 37826 47172 37832 47184
rect 35023 47144 37832 47172
rect 35023 47141 35035 47144
rect 34977 47135 35035 47141
rect 12989 47107 13047 47113
rect 12989 47073 13001 47107
rect 13035 47104 13047 47107
rect 13538 47104 13544 47116
rect 13035 47076 13544 47104
rect 13035 47073 13047 47076
rect 12989 47067 13047 47073
rect 13538 47064 13544 47076
rect 13596 47064 13602 47116
rect 14921 47107 14979 47113
rect 14921 47073 14933 47107
rect 14967 47104 14979 47107
rect 15562 47104 15568 47116
rect 14967 47076 15568 47104
rect 14967 47073 14979 47076
rect 14921 47067 14979 47073
rect 15562 47064 15568 47076
rect 15620 47064 15626 47116
rect 16298 47104 16304 47116
rect 16259 47076 16304 47104
rect 16298 47064 16304 47076
rect 16356 47064 16362 47116
rect 20162 47064 20168 47116
rect 20220 47104 20226 47116
rect 22097 47107 22155 47113
rect 22097 47104 22109 47107
rect 20220 47076 22109 47104
rect 20220 47064 20226 47076
rect 22097 47073 22109 47076
rect 22143 47073 22155 47107
rect 26418 47104 26424 47116
rect 26379 47076 26424 47104
rect 22097 47067 22155 47073
rect 26418 47064 26424 47076
rect 26476 47064 26482 47116
rect 29270 47064 29276 47116
rect 29328 47104 29334 47116
rect 33594 47104 33600 47116
rect 29328 47076 33600 47104
rect 29328 47064 29334 47076
rect 33594 47064 33600 47076
rect 33652 47064 33658 47116
rect 34330 47064 34336 47116
rect 34388 47104 34394 47116
rect 34992 47104 35020 47135
rect 37826 47132 37832 47144
rect 37884 47132 37890 47184
rect 34388 47076 35020 47104
rect 34388 47064 34394 47076
rect 35434 47064 35440 47116
rect 35492 47104 35498 47116
rect 35492 47076 35756 47104
rect 35492 47064 35498 47076
rect 2314 47036 2320 47048
rect 2275 47008 2320 47036
rect 2314 46996 2320 47008
rect 2372 47036 2378 47048
rect 6822 47036 6828 47048
rect 2372 47008 6828 47036
rect 2372 46996 2378 47008
rect 6822 46996 6828 47008
rect 6880 46996 6886 47048
rect 12345 47039 12403 47045
rect 12345 47005 12357 47039
rect 12391 47036 12403 47039
rect 12618 47036 12624 47048
rect 12391 47008 12624 47036
rect 12391 47005 12403 47008
rect 12345 46999 12403 47005
rect 12618 46996 12624 47008
rect 12676 46996 12682 47048
rect 13173 47039 13231 47045
rect 13173 47005 13185 47039
rect 13219 47036 13231 47039
rect 13262 47036 13268 47048
rect 13219 47008 13268 47036
rect 13219 47005 13231 47008
rect 13173 46999 13231 47005
rect 13262 46996 13268 47008
rect 13320 46996 13326 47048
rect 15105 47039 15163 47045
rect 15105 47005 15117 47039
rect 15151 47036 15163 47039
rect 15286 47036 15292 47048
rect 15151 47008 15292 47036
rect 15151 47005 15163 47008
rect 15105 46999 15163 47005
rect 15286 46996 15292 47008
rect 15344 46996 15350 47048
rect 16568 47039 16626 47045
rect 16568 47005 16580 47039
rect 16614 47036 16626 47039
rect 17034 47036 17040 47048
rect 16614 47008 17040 47036
rect 16614 47005 16626 47008
rect 16568 46999 16626 47005
rect 17034 46996 17040 47008
rect 17092 46996 17098 47048
rect 20257 47039 20315 47045
rect 20257 47005 20269 47039
rect 20303 47036 20315 47039
rect 20806 47036 20812 47048
rect 20303 47008 20812 47036
rect 20303 47005 20315 47008
rect 20257 46999 20315 47005
rect 20806 46996 20812 47008
rect 20864 46996 20870 47048
rect 20990 47036 20996 47048
rect 20951 47008 20996 47036
rect 20990 46996 20996 47008
rect 21048 46996 21054 47048
rect 21818 47036 21824 47048
rect 21731 47008 21824 47036
rect 21818 46996 21824 47008
rect 21876 46996 21882 47048
rect 23290 47036 23296 47048
rect 23251 47008 23296 47036
rect 23290 46996 23296 47008
rect 23348 46996 23354 47048
rect 26688 47039 26746 47045
rect 26688 47005 26700 47039
rect 26734 47036 26746 47039
rect 27154 47036 27160 47048
rect 26734 47008 27160 47036
rect 26734 47005 26746 47008
rect 26688 46999 26746 47005
rect 27154 46996 27160 47008
rect 27212 46996 27218 47048
rect 28721 47039 28779 47045
rect 28721 47005 28733 47039
rect 28767 47036 28779 47039
rect 29288 47036 29316 47064
rect 28767 47008 29316 47036
rect 28767 47005 28779 47008
rect 28721 46999 28779 47005
rect 31570 46996 31576 47048
rect 31628 47036 31634 47048
rect 31665 47039 31723 47045
rect 31665 47036 31677 47039
rect 31628 47008 31677 47036
rect 31628 46996 31634 47008
rect 31665 47005 31677 47008
rect 31711 47005 31723 47039
rect 32490 47036 32496 47048
rect 32451 47008 32496 47036
rect 31665 46999 31723 47005
rect 32490 46996 32496 47008
rect 32548 46996 32554 47048
rect 33612 47036 33640 47064
rect 35728 47045 35756 47076
rect 35802 47064 35808 47116
rect 35860 47104 35866 47116
rect 35860 47076 37504 47104
rect 35860 47064 35866 47076
rect 36096 47045 36124 47076
rect 35713 47039 35771 47045
rect 33612 47008 35664 47036
rect 21836 46968 21864 46996
rect 25590 46968 25596 46980
rect 21836 46940 25596 46968
rect 25590 46928 25596 46940
rect 25648 46928 25654 46980
rect 30190 46968 30196 46980
rect 30151 46940 30196 46968
rect 30190 46928 30196 46940
rect 30248 46928 30254 46980
rect 30282 46928 30288 46980
rect 30340 46968 30346 46980
rect 30393 46971 30451 46977
rect 30393 46968 30405 46971
rect 30340 46940 30405 46968
rect 30340 46928 30346 46940
rect 30393 46937 30405 46940
rect 30439 46937 30451 46971
rect 30393 46931 30451 46937
rect 30558 46928 30564 46980
rect 30616 46968 30622 46980
rect 33502 46968 33508 46980
rect 30616 46940 33508 46968
rect 30616 46928 30622 46940
rect 33502 46928 33508 46940
rect 33560 46928 33566 46980
rect 33778 46968 33784 46980
rect 33739 46940 33784 46968
rect 33778 46928 33784 46940
rect 33836 46928 33842 46980
rect 33997 46971 34055 46977
rect 33997 46937 34009 46971
rect 34043 46968 34055 46971
rect 34793 46971 34851 46977
rect 34793 46968 34805 46971
rect 34043 46940 34805 46968
rect 34043 46937 34055 46940
rect 33997 46931 34055 46937
rect 34793 46937 34805 46940
rect 34839 46968 34851 46971
rect 35526 46968 35532 46980
rect 34839 46940 35532 46968
rect 34839 46937 34851 46940
rect 34793 46931 34851 46937
rect 35526 46928 35532 46940
rect 35584 46928 35590 46980
rect 35636 46968 35664 47008
rect 35713 47005 35725 47039
rect 35759 47005 35771 47039
rect 35713 46999 35771 47005
rect 36081 47039 36139 47045
rect 36081 47005 36093 47039
rect 36127 47005 36139 47039
rect 36446 47036 36452 47048
rect 36407 47008 36452 47036
rect 36081 46999 36139 47005
rect 36446 46996 36452 47008
rect 36504 46996 36510 47048
rect 36722 47036 36728 47048
rect 36683 47008 36728 47036
rect 36722 46996 36728 47008
rect 36780 46996 36786 47048
rect 36354 46968 36360 46980
rect 35636 46940 36360 46968
rect 36354 46928 36360 46940
rect 36412 46928 36418 46980
rect 36633 46971 36691 46977
rect 36633 46937 36645 46971
rect 36679 46968 36691 46971
rect 37274 46968 37280 46980
rect 36679 46940 37280 46968
rect 36679 46937 36691 46940
rect 36633 46931 36691 46937
rect 37274 46928 37280 46940
rect 37332 46928 37338 46980
rect 19978 46860 19984 46912
rect 20036 46900 20042 46912
rect 20257 46903 20315 46909
rect 20257 46900 20269 46903
rect 20036 46872 20269 46900
rect 20036 46860 20042 46872
rect 20257 46869 20269 46872
rect 20303 46869 20315 46903
rect 20806 46900 20812 46912
rect 20767 46872 20812 46900
rect 20257 46863 20315 46869
rect 20806 46860 20812 46872
rect 20864 46860 20870 46912
rect 24026 46860 24032 46912
rect 24084 46900 24090 46912
rect 24854 46900 24860 46912
rect 24084 46872 24860 46900
rect 24084 46860 24090 46872
rect 24854 46860 24860 46872
rect 24912 46860 24918 46912
rect 28902 46900 28908 46912
rect 28863 46872 28908 46900
rect 28902 46860 28908 46872
rect 28960 46860 28966 46912
rect 31846 46900 31852 46912
rect 31807 46872 31852 46900
rect 31846 46860 31852 46872
rect 31904 46860 31910 46912
rect 32030 46860 32036 46912
rect 32088 46900 32094 46912
rect 37476 46909 37504 47076
rect 37645 47039 37703 47045
rect 37645 47005 37657 47039
rect 37691 47005 37703 47039
rect 38010 47036 38016 47048
rect 37971 47008 38016 47036
rect 37645 46999 37703 47005
rect 37660 46968 37688 46999
rect 38010 46996 38016 47008
rect 38068 46996 38074 47048
rect 38102 46996 38108 47048
rect 38160 47036 38166 47048
rect 38197 47039 38255 47045
rect 38197 47036 38209 47039
rect 38160 47008 38209 47036
rect 38160 46996 38166 47008
rect 38197 47005 38209 47008
rect 38243 47005 38255 47039
rect 38930 47036 38936 47048
rect 38891 47008 38936 47036
rect 38197 46999 38255 47005
rect 38930 46996 38936 47008
rect 38988 46996 38994 47048
rect 40052 47036 40080 47203
rect 40218 47200 40224 47212
rect 40276 47200 40282 47252
rect 44358 47200 44364 47252
rect 44416 47240 44422 47252
rect 45373 47243 45431 47249
rect 45373 47240 45385 47243
rect 44416 47212 45385 47240
rect 44416 47200 44422 47212
rect 45373 47209 45385 47212
rect 45419 47209 45431 47243
rect 45373 47203 45431 47209
rect 45833 47243 45891 47249
rect 45833 47209 45845 47243
rect 45879 47240 45891 47243
rect 46106 47240 46112 47252
rect 45879 47212 46112 47240
rect 45879 47209 45891 47212
rect 45833 47203 45891 47209
rect 46106 47200 46112 47212
rect 46164 47200 46170 47252
rect 46290 47240 46296 47252
rect 46251 47212 46296 47240
rect 46290 47200 46296 47212
rect 46348 47200 46354 47252
rect 46658 47240 46664 47252
rect 46619 47212 46664 47240
rect 46658 47200 46664 47212
rect 46716 47200 46722 47252
rect 51442 47200 51448 47252
rect 51500 47240 51506 47252
rect 53009 47243 53067 47249
rect 53009 47240 53021 47243
rect 51500 47212 53021 47240
rect 51500 47200 51506 47212
rect 53009 47209 53021 47212
rect 53055 47209 53067 47243
rect 53009 47203 53067 47209
rect 41233 47175 41291 47181
rect 41233 47141 41245 47175
rect 41279 47172 41291 47175
rect 41690 47172 41696 47184
rect 41279 47144 41696 47172
rect 41279 47141 41291 47144
rect 41233 47135 41291 47141
rect 41690 47132 41696 47144
rect 41748 47132 41754 47184
rect 40126 47064 40132 47116
rect 40184 47104 40190 47116
rect 40773 47107 40831 47113
rect 40773 47104 40785 47107
rect 40184 47076 40785 47104
rect 40184 47064 40190 47076
rect 40773 47073 40785 47076
rect 40819 47104 40831 47107
rect 40954 47104 40960 47116
rect 40819 47076 40960 47104
rect 40819 47073 40831 47076
rect 40773 47067 40831 47073
rect 40954 47064 40960 47076
rect 41012 47064 41018 47116
rect 45557 47107 45615 47113
rect 45557 47073 45569 47107
rect 45603 47104 45615 47107
rect 45830 47104 45836 47116
rect 45603 47076 45836 47104
rect 45603 47073 45615 47076
rect 45557 47067 45615 47073
rect 45830 47064 45836 47076
rect 45888 47064 45894 47116
rect 66990 47064 66996 47116
rect 67048 47104 67054 47116
rect 67174 47104 67180 47116
rect 67048 47076 67180 47104
rect 67048 47064 67054 47076
rect 67174 47064 67180 47076
rect 67232 47064 67238 47116
rect 40865 47039 40923 47045
rect 40865 47036 40877 47039
rect 40052 47008 40877 47036
rect 40865 47005 40877 47008
rect 40911 47036 40923 47039
rect 44177 47039 44235 47045
rect 44177 47036 44189 47039
rect 40911 47008 44189 47036
rect 40911 47005 40923 47008
rect 40865 46999 40923 47005
rect 44177 47005 44189 47008
rect 44223 47036 44235 47039
rect 44450 47036 44456 47048
rect 44223 47008 44456 47036
rect 44223 47005 44235 47008
rect 44177 46999 44235 47005
rect 44450 46996 44456 47008
rect 44508 46996 44514 47048
rect 44910 46996 44916 47048
rect 44968 47036 44974 47048
rect 45373 47039 45431 47045
rect 45373 47036 45385 47039
rect 44968 47008 45385 47036
rect 44968 46996 44974 47008
rect 45373 47005 45385 47008
rect 45419 47005 45431 47039
rect 45646 47036 45652 47048
rect 45607 47008 45652 47036
rect 45373 46999 45431 47005
rect 37918 46968 37924 46980
rect 37660 46940 37924 46968
rect 37918 46928 37924 46940
rect 37976 46928 37982 46980
rect 39853 46971 39911 46977
rect 39853 46937 39865 46971
rect 39899 46968 39911 46971
rect 39942 46968 39948 46980
rect 39899 46940 39948 46968
rect 39899 46937 39911 46940
rect 39853 46931 39911 46937
rect 39942 46928 39948 46940
rect 40000 46928 40006 46980
rect 40034 46928 40040 46980
rect 40092 46977 40098 46980
rect 40092 46971 40111 46977
rect 40099 46937 40111 46971
rect 40092 46931 40111 46937
rect 40092 46928 40098 46931
rect 43438 46928 43444 46980
rect 43496 46968 43502 46980
rect 43993 46971 44051 46977
rect 43993 46968 44005 46971
rect 43496 46940 44005 46968
rect 43496 46928 43502 46940
rect 43993 46937 44005 46940
rect 44039 46968 44051 46971
rect 45388 46968 45416 46999
rect 45646 46996 45652 47008
rect 45704 46996 45710 47048
rect 46293 47039 46351 47045
rect 46293 47005 46305 47039
rect 46339 47005 46351 47039
rect 46293 46999 46351 47005
rect 46308 46968 46336 46999
rect 46382 46996 46388 47048
rect 46440 47036 46446 47048
rect 50985 47039 51043 47045
rect 46440 47008 46485 47036
rect 46440 46996 46446 47008
rect 50985 47005 50997 47039
rect 51031 47005 51043 47039
rect 50985 46999 51043 47005
rect 51169 47039 51227 47045
rect 51169 47005 51181 47039
rect 51215 47036 51227 47039
rect 51629 47039 51687 47045
rect 51629 47036 51641 47039
rect 51215 47008 51641 47036
rect 51215 47005 51227 47008
rect 51169 46999 51227 47005
rect 51629 47005 51641 47008
rect 51675 47005 51687 47039
rect 51629 46999 51687 47005
rect 44039 46940 44220 46968
rect 45388 46940 46336 46968
rect 51000 46968 51028 46999
rect 51718 46996 51724 47048
rect 51776 47036 51782 47048
rect 51885 47039 51943 47045
rect 51885 47036 51897 47039
rect 51776 47008 51897 47036
rect 51776 46996 51782 47008
rect 51885 47005 51897 47008
rect 51931 47005 51943 47039
rect 51885 46999 51943 47005
rect 66254 46996 66260 47048
rect 66312 47036 66318 47048
rect 67913 47039 67971 47045
rect 67913 47036 67925 47039
rect 66312 47008 67925 47036
rect 66312 46996 66318 47008
rect 67913 47005 67925 47008
rect 67959 47005 67971 47039
rect 67913 46999 67971 47005
rect 51350 46968 51356 46980
rect 51000 46940 51356 46968
rect 44039 46937 44051 46940
rect 43993 46931 44051 46937
rect 32585 46903 32643 46909
rect 32585 46900 32597 46903
rect 32088 46872 32597 46900
rect 32088 46860 32094 46872
rect 32585 46869 32597 46872
rect 32631 46869 32643 46903
rect 32585 46863 32643 46869
rect 37461 46903 37519 46909
rect 37461 46869 37473 46903
rect 37507 46869 37519 46903
rect 44192 46900 44220 46940
rect 51350 46928 51356 46940
rect 51408 46928 51414 46980
rect 58710 46928 58716 46980
rect 58768 46968 58774 46980
rect 67082 46968 67088 46980
rect 58768 46940 67088 46968
rect 58768 46928 58774 46940
rect 67082 46928 67088 46940
rect 67140 46928 67146 46980
rect 46382 46900 46388 46912
rect 44192 46872 46388 46900
rect 37461 46863 37519 46869
rect 46382 46860 46388 46872
rect 46440 46860 46446 46912
rect 1104 46810 68816 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 68816 46810
rect 1104 46736 68816 46758
rect 22094 46656 22100 46708
rect 22152 46696 22158 46708
rect 22152 46668 26234 46696
rect 22152 46656 22158 46668
rect 17310 46588 17316 46640
rect 17368 46628 17374 46640
rect 20156 46631 20214 46637
rect 17368 46600 17540 46628
rect 17368 46588 17374 46600
rect 17512 46572 17540 46600
rect 20156 46597 20168 46631
rect 20202 46628 20214 46631
rect 20806 46628 20812 46640
rect 20202 46600 20812 46628
rect 20202 46597 20214 46600
rect 20156 46591 20214 46597
rect 20806 46588 20812 46600
rect 20864 46588 20870 46640
rect 26206 46628 26234 46668
rect 28626 46656 28632 46708
rect 28684 46696 28690 46708
rect 32950 46696 32956 46708
rect 28684 46668 32956 46696
rect 28684 46656 28690 46668
rect 32950 46656 32956 46668
rect 33008 46656 33014 46708
rect 35618 46656 35624 46708
rect 35676 46696 35682 46708
rect 36262 46696 36268 46708
rect 35676 46668 36268 46696
rect 35676 46656 35682 46668
rect 36262 46656 36268 46668
rect 36320 46696 36326 46708
rect 36449 46699 36507 46705
rect 36449 46696 36461 46699
rect 36320 46668 36461 46696
rect 36320 46656 36326 46668
rect 36449 46665 36461 46668
rect 36495 46665 36507 46699
rect 42610 46696 42616 46708
rect 42571 46668 42616 46696
rect 36449 46659 36507 46665
rect 42610 46656 42616 46668
rect 42668 46656 42674 46708
rect 43162 46696 43168 46708
rect 43123 46668 43168 46696
rect 43162 46656 43168 46668
rect 43220 46656 43226 46708
rect 45554 46656 45560 46708
rect 45612 46696 45618 46708
rect 45833 46699 45891 46705
rect 45833 46696 45845 46699
rect 45612 46668 45845 46696
rect 45612 46656 45618 46668
rect 45833 46665 45845 46668
rect 45879 46665 45891 46699
rect 45833 46659 45891 46665
rect 47578 46656 47584 46708
rect 47636 46696 47642 46708
rect 48961 46699 49019 46705
rect 48961 46696 48973 46699
rect 47636 46668 48973 46696
rect 47636 46656 47642 46668
rect 48961 46665 48973 46668
rect 49007 46665 49019 46699
rect 50798 46696 50804 46708
rect 50759 46668 50804 46696
rect 48961 46659 49019 46665
rect 50798 46656 50804 46668
rect 50856 46656 50862 46708
rect 51626 46656 51632 46708
rect 51684 46696 51690 46708
rect 51905 46699 51963 46705
rect 51905 46696 51917 46699
rect 51684 46668 51917 46696
rect 51684 46656 51690 46668
rect 51905 46665 51917 46668
rect 51951 46665 51963 46699
rect 51905 46659 51963 46665
rect 34057 46631 34115 46637
rect 34057 46628 34069 46631
rect 26206 46600 34069 46628
rect 34057 46597 34069 46600
rect 34103 46597 34115 46631
rect 40218 46628 40224 46640
rect 34057 46591 34115 46597
rect 39408 46600 40224 46628
rect 1854 46560 1860 46572
rect 1815 46532 1860 46560
rect 1854 46520 1860 46532
rect 1912 46520 1918 46572
rect 17402 46560 17408 46572
rect 17363 46532 17408 46560
rect 17402 46520 17408 46532
rect 17460 46520 17466 46572
rect 17494 46520 17500 46572
rect 17552 46560 17558 46572
rect 17552 46532 17645 46560
rect 17552 46520 17558 46532
rect 18966 46520 18972 46572
rect 19024 46560 19030 46572
rect 19061 46563 19119 46569
rect 19061 46560 19073 46563
rect 19024 46532 19073 46560
rect 19024 46520 19030 46532
rect 19061 46529 19073 46532
rect 19107 46529 19119 46563
rect 19061 46523 19119 46529
rect 19889 46563 19947 46569
rect 19889 46529 19901 46563
rect 19935 46560 19947 46563
rect 19978 46560 19984 46572
rect 19935 46532 19984 46560
rect 19935 46529 19947 46532
rect 19889 46523 19947 46529
rect 19978 46520 19984 46532
rect 20036 46520 20042 46572
rect 20898 46520 20904 46572
rect 20956 46560 20962 46572
rect 21821 46563 21879 46569
rect 21821 46560 21833 46563
rect 20956 46532 21833 46560
rect 20956 46520 20962 46532
rect 21821 46529 21833 46532
rect 21867 46529 21879 46563
rect 21821 46523 21879 46529
rect 22278 46520 22284 46572
rect 22336 46560 22342 46572
rect 22741 46563 22799 46569
rect 22741 46560 22753 46563
rect 22336 46532 22753 46560
rect 22336 46520 22342 46532
rect 22741 46529 22753 46532
rect 22787 46529 22799 46563
rect 24026 46560 24032 46572
rect 23987 46532 24032 46560
rect 22741 46523 22799 46529
rect 24026 46520 24032 46532
rect 24084 46520 24090 46572
rect 24946 46520 24952 46572
rect 25004 46560 25010 46572
rect 25004 46532 25049 46560
rect 25004 46520 25010 46532
rect 27982 46520 27988 46572
rect 28040 46560 28046 46572
rect 28537 46563 28595 46569
rect 28537 46560 28549 46563
rect 28040 46532 28549 46560
rect 28040 46520 28046 46532
rect 28537 46529 28549 46532
rect 28583 46560 28595 46563
rect 28902 46560 28908 46572
rect 28583 46532 28908 46560
rect 28583 46529 28595 46532
rect 28537 46523 28595 46529
rect 28902 46520 28908 46532
rect 28960 46520 28966 46572
rect 29270 46560 29276 46572
rect 29231 46532 29276 46560
rect 29270 46520 29276 46532
rect 29328 46520 29334 46572
rect 30006 46560 30012 46572
rect 29967 46532 30012 46560
rect 30006 46520 30012 46532
rect 30064 46520 30070 46572
rect 30926 46560 30932 46572
rect 30887 46532 30932 46560
rect 30926 46520 30932 46532
rect 30984 46520 30990 46572
rect 33410 46560 33416 46572
rect 32784 46532 33416 46560
rect 24213 46495 24271 46501
rect 24213 46461 24225 46495
rect 24259 46492 24271 46495
rect 24762 46492 24768 46504
rect 24259 46464 24768 46492
rect 24259 46461 24271 46464
rect 24213 46455 24271 46461
rect 24762 46452 24768 46464
rect 24820 46452 24826 46504
rect 25038 46452 25044 46504
rect 25096 46501 25102 46504
rect 25096 46495 25124 46501
rect 25112 46461 25124 46495
rect 25096 46455 25124 46461
rect 25225 46495 25283 46501
rect 25225 46461 25237 46495
rect 25271 46492 25283 46495
rect 26050 46492 26056 46504
rect 25271 46464 26056 46492
rect 25271 46461 25283 46464
rect 25225 46455 25283 46461
rect 25096 46452 25102 46455
rect 26050 46452 26056 46464
rect 26108 46452 26114 46504
rect 30024 46492 30052 46520
rect 32784 46504 32812 46532
rect 33410 46520 33416 46532
rect 33468 46520 33474 46572
rect 35894 46520 35900 46572
rect 35952 46560 35958 46572
rect 36357 46563 36415 46569
rect 36357 46560 36369 46563
rect 35952 46532 36369 46560
rect 35952 46520 35958 46532
rect 36357 46529 36369 46532
rect 36403 46560 36415 46563
rect 36722 46560 36728 46572
rect 36403 46532 36728 46560
rect 36403 46529 36415 46532
rect 36357 46523 36415 46529
rect 36722 46520 36728 46532
rect 36780 46520 36786 46572
rect 37274 46520 37280 46572
rect 37332 46560 37338 46572
rect 37737 46563 37795 46569
rect 37737 46560 37749 46563
rect 37332 46532 37749 46560
rect 37332 46520 37338 46532
rect 37737 46529 37749 46532
rect 37783 46560 37795 46563
rect 38562 46560 38568 46572
rect 37783 46532 38568 46560
rect 37783 46529 37795 46532
rect 37737 46523 37795 46529
rect 38562 46520 38568 46532
rect 38620 46520 38626 46572
rect 39408 46569 39436 46600
rect 40218 46588 40224 46600
rect 40276 46588 40282 46640
rect 42058 46628 42064 46640
rect 41892 46600 42064 46628
rect 39393 46563 39451 46569
rect 39393 46529 39405 46563
rect 39439 46529 39451 46563
rect 39393 46523 39451 46529
rect 39485 46563 39543 46569
rect 39485 46529 39497 46563
rect 39531 46560 39543 46563
rect 40678 46560 40684 46572
rect 39531 46532 40684 46560
rect 39531 46529 39543 46532
rect 39485 46523 39543 46529
rect 40678 46520 40684 46532
rect 40736 46520 40742 46572
rect 41690 46560 41696 46572
rect 41651 46532 41696 46560
rect 41690 46520 41696 46532
rect 41748 46520 41754 46572
rect 41892 46569 41920 46600
rect 42058 46588 42064 46600
rect 42116 46628 42122 46640
rect 47118 46628 47124 46640
rect 42116 46600 47124 46628
rect 42116 46588 42122 46600
rect 47118 46588 47124 46600
rect 47176 46588 47182 46640
rect 47210 46588 47216 46640
rect 47268 46628 47274 46640
rect 47826 46631 47884 46637
rect 47826 46628 47838 46631
rect 47268 46600 47838 46628
rect 47268 46588 47274 46600
rect 47826 46597 47838 46600
rect 47872 46597 47884 46631
rect 47826 46591 47884 46597
rect 48038 46588 48044 46640
rect 48096 46588 48102 46640
rect 49694 46637 49700 46640
rect 49688 46628 49700 46637
rect 49655 46600 49700 46628
rect 49688 46591 49700 46600
rect 49694 46588 49700 46591
rect 49752 46588 49758 46640
rect 66254 46628 66260 46640
rect 65812 46600 66260 46628
rect 41877 46563 41935 46569
rect 41877 46529 41889 46563
rect 41923 46529 41935 46563
rect 41877 46523 41935 46529
rect 42426 46520 42432 46572
rect 42484 46560 42490 46572
rect 42521 46563 42579 46569
rect 42521 46560 42533 46563
rect 42484 46532 42533 46560
rect 42484 46520 42490 46532
rect 42521 46529 42533 46532
rect 42567 46560 42579 46563
rect 43349 46563 43407 46569
rect 43349 46560 43361 46563
rect 42567 46532 43361 46560
rect 42567 46529 42579 46532
rect 42521 46523 42579 46529
rect 43349 46529 43361 46532
rect 43395 46529 43407 46563
rect 43349 46523 43407 46529
rect 43625 46563 43683 46569
rect 43625 46529 43637 46563
rect 43671 46560 43683 46563
rect 43898 46560 43904 46572
rect 43671 46532 43904 46560
rect 43671 46529 43683 46532
rect 43625 46523 43683 46529
rect 43898 46520 43904 46532
rect 43956 46520 43962 46572
rect 44358 46520 44364 46572
rect 44416 46560 44422 46572
rect 44453 46563 44511 46569
rect 44453 46560 44465 46563
rect 44416 46532 44465 46560
rect 44416 46520 44422 46532
rect 44453 46529 44465 46532
rect 44499 46529 44511 46563
rect 44453 46523 44511 46529
rect 45465 46563 45523 46569
rect 45465 46529 45477 46563
rect 45511 46529 45523 46563
rect 45646 46560 45652 46572
rect 45607 46532 45652 46560
rect 45465 46523 45523 46529
rect 31846 46492 31852 46504
rect 30024 46464 31852 46492
rect 31846 46452 31852 46464
rect 31904 46492 31910 46504
rect 32490 46492 32496 46504
rect 31904 46464 32496 46492
rect 31904 46452 31910 46464
rect 32490 46452 32496 46464
rect 32548 46452 32554 46504
rect 32766 46492 32772 46504
rect 32727 46464 32772 46492
rect 32766 46452 32772 46464
rect 32824 46452 32830 46504
rect 32858 46452 32864 46504
rect 32916 46492 32922 46504
rect 33045 46495 33103 46501
rect 33045 46492 33057 46495
rect 32916 46464 33057 46492
rect 32916 46452 32922 46464
rect 33045 46461 33057 46464
rect 33091 46461 33103 46495
rect 33045 46455 33103 46461
rect 35342 46452 35348 46504
rect 35400 46492 35406 46504
rect 35805 46495 35863 46501
rect 35805 46492 35817 46495
rect 35400 46464 35817 46492
rect 35400 46452 35406 46464
rect 35805 46461 35817 46464
rect 35851 46492 35863 46495
rect 38194 46492 38200 46504
rect 35851 46464 38200 46492
rect 35851 46461 35863 46464
rect 35805 46455 35863 46461
rect 38194 46452 38200 46464
rect 38252 46452 38258 46504
rect 39669 46495 39727 46501
rect 39669 46461 39681 46495
rect 39715 46492 39727 46495
rect 39942 46492 39948 46504
rect 39715 46464 39948 46492
rect 39715 46461 39727 46464
rect 39669 46455 39727 46461
rect 39942 46452 39948 46464
rect 40000 46452 40006 46504
rect 44177 46495 44235 46501
rect 44177 46461 44189 46495
rect 44223 46461 44235 46495
rect 44177 46455 44235 46461
rect 2038 46424 2044 46436
rect 1999 46396 2044 46424
rect 2038 46384 2044 46396
rect 2096 46384 2102 46436
rect 24673 46427 24731 46433
rect 24673 46393 24685 46427
rect 24719 46393 24731 46427
rect 24673 46387 24731 46393
rect 25608 46396 26234 46424
rect 17681 46359 17739 46365
rect 17681 46325 17693 46359
rect 17727 46356 17739 46359
rect 18506 46356 18512 46368
rect 17727 46328 18512 46356
rect 17727 46325 17739 46328
rect 17681 46319 17739 46325
rect 18506 46316 18512 46328
rect 18564 46316 18570 46368
rect 19242 46356 19248 46368
rect 19203 46328 19248 46356
rect 19242 46316 19248 46328
rect 19300 46316 19306 46368
rect 19702 46316 19708 46368
rect 19760 46356 19766 46368
rect 21269 46359 21327 46365
rect 21269 46356 21281 46359
rect 19760 46328 21281 46356
rect 19760 46316 19766 46328
rect 21269 46325 21281 46328
rect 21315 46325 21327 46359
rect 21269 46319 21327 46325
rect 21634 46316 21640 46368
rect 21692 46356 21698 46368
rect 21821 46359 21879 46365
rect 21821 46356 21833 46359
rect 21692 46328 21833 46356
rect 21692 46316 21698 46328
rect 21821 46325 21833 46328
rect 21867 46325 21879 46359
rect 21821 46319 21879 46325
rect 21910 46316 21916 46368
rect 21968 46356 21974 46368
rect 22557 46359 22615 46365
rect 22557 46356 22569 46359
rect 21968 46328 22569 46356
rect 21968 46316 21974 46328
rect 22557 46325 22569 46328
rect 22603 46325 22615 46359
rect 24688 46356 24716 46387
rect 25608 46356 25636 46396
rect 24688 46328 25636 46356
rect 22557 46319 22615 46325
rect 25682 46316 25688 46368
rect 25740 46356 25746 46368
rect 25869 46359 25927 46365
rect 25869 46356 25881 46359
rect 25740 46328 25881 46356
rect 25740 46316 25746 46328
rect 25869 46325 25881 46328
rect 25915 46325 25927 46359
rect 26206 46356 26234 46396
rect 26326 46384 26332 46436
rect 26384 46424 26390 46436
rect 33778 46424 33784 46436
rect 26384 46396 33784 46424
rect 26384 46384 26390 46396
rect 33778 46384 33784 46396
rect 33836 46384 33842 46436
rect 38013 46427 38071 46433
rect 38013 46393 38025 46427
rect 38059 46424 38071 46427
rect 38286 46424 38292 46436
rect 38059 46396 38292 46424
rect 38059 46393 38071 46396
rect 38013 46387 38071 46393
rect 38286 46384 38292 46396
rect 38344 46424 38350 46436
rect 39022 46424 39028 46436
rect 38344 46396 39028 46424
rect 38344 46384 38350 46396
rect 39022 46384 39028 46396
rect 39080 46384 39086 46436
rect 43438 46424 43444 46436
rect 43399 46396 43444 46424
rect 43438 46384 43444 46396
rect 43496 46384 43502 46436
rect 43530 46384 43536 46436
rect 43588 46424 43594 46436
rect 44192 46424 44220 46455
rect 43588 46396 44220 46424
rect 43588 46384 43594 46396
rect 28626 46356 28632 46368
rect 26206 46328 28632 46356
rect 25869 46319 25927 46325
rect 28626 46316 28632 46328
rect 28684 46316 28690 46368
rect 28994 46316 29000 46368
rect 29052 46356 29058 46368
rect 29362 46356 29368 46368
rect 29052 46328 29368 46356
rect 29052 46316 29058 46328
rect 29362 46316 29368 46328
rect 29420 46356 29426 46368
rect 29457 46359 29515 46365
rect 29457 46356 29469 46359
rect 29420 46328 29469 46356
rect 29420 46316 29426 46328
rect 29457 46325 29469 46328
rect 29503 46325 29515 46359
rect 29457 46319 29515 46325
rect 29914 46316 29920 46368
rect 29972 46356 29978 46368
rect 30009 46359 30067 46365
rect 30009 46356 30021 46359
rect 29972 46328 30021 46356
rect 29972 46316 29978 46328
rect 30009 46325 30021 46328
rect 30055 46325 30067 46359
rect 30742 46356 30748 46368
rect 30703 46328 30748 46356
rect 30009 46319 30067 46325
rect 30742 46316 30748 46328
rect 30800 46316 30806 46368
rect 38654 46316 38660 46368
rect 38712 46356 38718 46368
rect 38749 46359 38807 46365
rect 38749 46356 38761 46359
rect 38712 46328 38761 46356
rect 38712 46316 38718 46328
rect 38749 46325 38761 46328
rect 38795 46356 38807 46359
rect 39114 46356 39120 46368
rect 38795 46328 39120 46356
rect 38795 46325 38807 46328
rect 38749 46319 38807 46325
rect 39114 46316 39120 46328
rect 39172 46316 39178 46368
rect 39577 46359 39635 46365
rect 39577 46325 39589 46359
rect 39623 46356 39635 46359
rect 40126 46356 40132 46368
rect 39623 46328 40132 46356
rect 39623 46325 39635 46328
rect 39577 46319 39635 46325
rect 40126 46316 40132 46328
rect 40184 46316 40190 46368
rect 41785 46359 41843 46365
rect 41785 46325 41797 46359
rect 41831 46356 41843 46359
rect 42150 46356 42156 46368
rect 41831 46328 42156 46356
rect 41831 46325 41843 46328
rect 41785 46319 41843 46325
rect 42150 46316 42156 46328
rect 42208 46316 42214 46368
rect 44468 46356 44496 46523
rect 45480 46492 45508 46523
rect 45646 46520 45652 46532
rect 45704 46520 45710 46572
rect 46937 46563 46995 46569
rect 46937 46529 46949 46563
rect 46983 46560 46995 46563
rect 48056 46560 48084 46588
rect 46983 46532 48084 46560
rect 46983 46529 46995 46532
rect 46937 46523 46995 46529
rect 51442 46520 51448 46572
rect 51500 46560 51506 46572
rect 51537 46563 51595 46569
rect 51537 46560 51549 46563
rect 51500 46532 51549 46560
rect 51500 46520 51506 46532
rect 51537 46529 51549 46532
rect 51583 46529 51595 46563
rect 51718 46560 51724 46572
rect 51679 46532 51724 46560
rect 51537 46523 51595 46529
rect 51718 46520 51724 46532
rect 51776 46520 51782 46572
rect 65812 46569 65840 46600
rect 66254 46588 66260 46600
rect 66312 46588 66318 46640
rect 65797 46563 65855 46569
rect 65797 46529 65809 46563
rect 65843 46529 65855 46563
rect 65797 46523 65855 46529
rect 45830 46492 45836 46504
rect 45480 46464 45836 46492
rect 45830 46452 45836 46464
rect 45888 46452 45894 46504
rect 47029 46495 47087 46501
rect 47029 46461 47041 46495
rect 47075 46492 47087 46495
rect 47581 46495 47639 46501
rect 47581 46492 47593 46495
rect 47075 46464 47593 46492
rect 47075 46461 47087 46464
rect 47029 46455 47087 46461
rect 47581 46461 47593 46464
rect 47627 46461 47639 46495
rect 49418 46492 49424 46504
rect 49379 46464 49424 46492
rect 47581 46455 47639 46461
rect 49418 46452 49424 46464
rect 49476 46452 49482 46504
rect 65981 46495 66039 46501
rect 65981 46461 65993 46495
rect 66027 46492 66039 46495
rect 67358 46492 67364 46504
rect 66027 46464 67364 46492
rect 66027 46461 66039 46464
rect 65981 46455 66039 46461
rect 67358 46452 67364 46464
rect 67416 46452 67422 46504
rect 67542 46492 67548 46504
rect 67503 46464 67548 46492
rect 67542 46452 67548 46464
rect 67600 46452 67606 46504
rect 45094 46356 45100 46368
rect 44468 46328 45100 46356
rect 45094 46316 45100 46328
rect 45152 46356 45158 46368
rect 45465 46359 45523 46365
rect 45465 46356 45477 46359
rect 45152 46328 45477 46356
rect 45152 46316 45158 46328
rect 45465 46325 45477 46328
rect 45511 46325 45523 46359
rect 45465 46319 45523 46325
rect 1104 46266 68816 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 65654 46266
rect 65706 46214 65718 46266
rect 65770 46214 65782 46266
rect 65834 46214 65846 46266
rect 65898 46214 65910 46266
rect 65962 46214 68816 46266
rect 1104 46192 68816 46214
rect 17402 46112 17408 46164
rect 17460 46152 17466 46164
rect 17865 46155 17923 46161
rect 17865 46152 17877 46155
rect 17460 46124 17877 46152
rect 17460 46112 17466 46124
rect 17865 46121 17877 46124
rect 17911 46121 17923 46155
rect 17865 46115 17923 46121
rect 19889 46155 19947 46161
rect 19889 46121 19901 46155
rect 19935 46152 19947 46155
rect 19978 46152 19984 46164
rect 19935 46124 19984 46152
rect 19935 46121 19947 46124
rect 19889 46115 19947 46121
rect 19978 46112 19984 46124
rect 20036 46152 20042 46164
rect 20717 46155 20775 46161
rect 20717 46152 20729 46155
rect 20036 46124 20729 46152
rect 20036 46112 20042 46124
rect 20717 46121 20729 46124
rect 20763 46121 20775 46155
rect 20717 46115 20775 46121
rect 21100 46124 22600 46152
rect 20073 46087 20131 46093
rect 20073 46053 20085 46087
rect 20119 46084 20131 46087
rect 20990 46084 20996 46096
rect 20119 46056 20996 46084
rect 20119 46053 20131 46056
rect 20073 46047 20131 46053
rect 20990 46044 20996 46056
rect 21048 46044 21054 46096
rect 19242 45976 19248 46028
rect 19300 46016 19306 46028
rect 21100 46016 21128 46124
rect 22572 46084 22600 46124
rect 24026 46112 24032 46164
rect 24084 46152 24090 46164
rect 25682 46152 25688 46164
rect 24084 46124 25688 46152
rect 24084 46112 24090 46124
rect 25682 46112 25688 46124
rect 25740 46112 25746 46164
rect 26050 46152 26056 46164
rect 25792 46124 26056 46152
rect 25792 46084 25820 46124
rect 26050 46112 26056 46124
rect 26108 46112 26114 46164
rect 33502 46112 33508 46164
rect 33560 46152 33566 46164
rect 35069 46155 35127 46161
rect 35069 46152 35081 46155
rect 33560 46124 35081 46152
rect 33560 46112 33566 46124
rect 35069 46121 35081 46124
rect 35115 46121 35127 46155
rect 35069 46115 35127 46121
rect 36170 46112 36176 46164
rect 36228 46152 36234 46164
rect 36817 46155 36875 46161
rect 36817 46152 36829 46155
rect 36228 46124 36829 46152
rect 36228 46112 36234 46124
rect 36817 46121 36829 46124
rect 36863 46121 36875 46155
rect 36817 46115 36875 46121
rect 41417 46155 41475 46161
rect 41417 46121 41429 46155
rect 41463 46152 41475 46155
rect 42426 46152 42432 46164
rect 41463 46124 42432 46152
rect 41463 46121 41475 46124
rect 41417 46115 41475 46121
rect 42426 46112 42432 46124
rect 42484 46112 42490 46164
rect 43438 46152 43444 46164
rect 43399 46124 43444 46152
rect 43438 46112 43444 46124
rect 43496 46112 43502 46164
rect 45189 46155 45247 46161
rect 45189 46121 45201 46155
rect 45235 46152 45247 46155
rect 45278 46152 45284 46164
rect 45235 46124 45284 46152
rect 45235 46121 45247 46124
rect 45189 46115 45247 46121
rect 45278 46112 45284 46124
rect 45336 46112 45342 46164
rect 45646 46112 45652 46164
rect 45704 46152 45710 46164
rect 45833 46155 45891 46161
rect 45833 46152 45845 46155
rect 45704 46124 45845 46152
rect 45704 46112 45710 46124
rect 45833 46121 45845 46124
rect 45879 46121 45891 46155
rect 45833 46115 45891 46121
rect 48225 46155 48283 46161
rect 48225 46121 48237 46155
rect 48271 46152 48283 46155
rect 49418 46152 49424 46164
rect 48271 46124 49424 46152
rect 48271 46121 48283 46124
rect 48225 46115 48283 46121
rect 49418 46112 49424 46124
rect 49476 46112 49482 46164
rect 66806 46112 66812 46164
rect 66864 46152 66870 46164
rect 67174 46152 67180 46164
rect 66864 46124 67180 46152
rect 66864 46112 66870 46124
rect 67174 46112 67180 46124
rect 67232 46112 67238 46164
rect 67358 46152 67364 46164
rect 67319 46124 67364 46152
rect 67358 46112 67364 46124
rect 67416 46112 67422 46164
rect 45094 46084 45100 46096
rect 22572 46056 25820 46084
rect 45055 46056 45100 46084
rect 45094 46044 45100 46056
rect 45152 46044 45158 46096
rect 21634 46016 21640 46028
rect 19300 45988 21128 46016
rect 21595 45988 21640 46016
rect 19300 45976 19306 45988
rect 21634 45976 21640 45988
rect 21692 45976 21698 46028
rect 24765 46019 24823 46025
rect 24765 46016 24777 46019
rect 23860 45988 24777 46016
rect 13173 45951 13231 45957
rect 13173 45917 13185 45951
rect 13219 45948 13231 45951
rect 13538 45948 13544 45960
rect 13219 45920 13544 45948
rect 13219 45917 13231 45920
rect 13173 45911 13231 45917
rect 13538 45908 13544 45920
rect 13596 45908 13602 45960
rect 14458 45948 14464 45960
rect 14419 45920 14464 45948
rect 14458 45908 14464 45920
rect 14516 45908 14522 45960
rect 15381 45951 15439 45957
rect 15381 45917 15393 45951
rect 15427 45948 15439 45951
rect 15470 45948 15476 45960
rect 15427 45920 15476 45948
rect 15427 45917 15439 45920
rect 15381 45911 15439 45917
rect 15470 45908 15476 45920
rect 15528 45908 15534 45960
rect 16485 45951 16543 45957
rect 16485 45917 16497 45951
rect 16531 45948 16543 45951
rect 16574 45948 16580 45960
rect 16531 45920 16580 45948
rect 16531 45917 16543 45920
rect 16485 45911 16543 45917
rect 16574 45908 16580 45920
rect 16632 45908 16638 45960
rect 18506 45948 18512 45960
rect 18467 45920 18512 45948
rect 18506 45908 18512 45920
rect 18564 45908 18570 45960
rect 18966 45908 18972 45960
rect 19024 45948 19030 45960
rect 21910 45957 21916 45960
rect 21904 45948 21916 45957
rect 19024 45920 20668 45948
rect 21871 45920 21916 45948
rect 19024 45908 19030 45920
rect 16752 45883 16810 45889
rect 16752 45849 16764 45883
rect 16798 45880 16810 45883
rect 16798 45852 18368 45880
rect 16798 45849 16810 45852
rect 16752 45843 16810 45849
rect 12986 45812 12992 45824
rect 12947 45784 12992 45812
rect 12986 45772 12992 45784
rect 13044 45772 13050 45824
rect 14642 45812 14648 45824
rect 14603 45784 14648 45812
rect 14642 45772 14648 45784
rect 14700 45772 14706 45824
rect 15194 45812 15200 45824
rect 15155 45784 15200 45812
rect 15194 45772 15200 45784
rect 15252 45772 15258 45824
rect 18340 45821 18368 45852
rect 19242 45840 19248 45892
rect 19300 45880 19306 45892
rect 19702 45880 19708 45892
rect 19300 45852 19708 45880
rect 19300 45840 19306 45852
rect 19702 45840 19708 45852
rect 19760 45840 19766 45892
rect 19921 45883 19979 45889
rect 19921 45849 19933 45883
rect 19967 45880 19979 45883
rect 20162 45880 20168 45892
rect 19967 45852 20168 45880
rect 19967 45849 19979 45852
rect 19921 45843 19979 45849
rect 20162 45840 20168 45852
rect 20220 45840 20226 45892
rect 20530 45880 20536 45892
rect 20491 45852 20536 45880
rect 20530 45840 20536 45852
rect 20588 45840 20594 45892
rect 20640 45880 20668 45920
rect 21904 45911 21916 45920
rect 21910 45908 21916 45911
rect 21968 45908 21974 45960
rect 23860 45957 23888 45988
rect 24765 45985 24777 45988
rect 24811 45985 24823 46019
rect 29914 46016 29920 46028
rect 24765 45979 24823 45985
rect 25148 45988 25912 46016
rect 29875 45988 29920 46016
rect 23845 45951 23903 45957
rect 23845 45917 23857 45951
rect 23891 45917 23903 45951
rect 23845 45911 23903 45917
rect 24489 45951 24547 45957
rect 24489 45917 24501 45951
rect 24535 45917 24547 45951
rect 24489 45911 24547 45917
rect 24581 45951 24639 45957
rect 24581 45917 24593 45951
rect 24627 45948 24639 45951
rect 24946 45948 24952 45960
rect 24627 45920 24952 45948
rect 24627 45917 24639 45920
rect 24581 45911 24639 45917
rect 24504 45880 24532 45911
rect 24946 45908 24952 45920
rect 25004 45908 25010 45960
rect 24670 45880 24676 45892
rect 20640 45852 23796 45880
rect 24504 45852 24676 45880
rect 18325 45815 18383 45821
rect 18325 45781 18337 45815
rect 18371 45781 18383 45815
rect 20180 45812 20208 45840
rect 20622 45812 20628 45824
rect 20180 45784 20628 45812
rect 18325 45775 18383 45781
rect 20622 45772 20628 45784
rect 20680 45812 20686 45824
rect 20733 45815 20791 45821
rect 20733 45812 20745 45815
rect 20680 45784 20745 45812
rect 20680 45772 20686 45784
rect 20733 45781 20745 45784
rect 20779 45781 20791 45815
rect 20898 45812 20904 45824
rect 20859 45784 20904 45812
rect 20733 45775 20791 45781
rect 20898 45772 20904 45784
rect 20956 45772 20962 45824
rect 21634 45772 21640 45824
rect 21692 45812 21698 45824
rect 23017 45815 23075 45821
rect 23017 45812 23029 45815
rect 21692 45784 23029 45812
rect 21692 45772 21698 45784
rect 23017 45781 23029 45784
rect 23063 45781 23075 45815
rect 23658 45812 23664 45824
rect 23619 45784 23664 45812
rect 23017 45775 23075 45781
rect 23658 45772 23664 45784
rect 23716 45772 23722 45824
rect 23768 45812 23796 45852
rect 24670 45840 24676 45852
rect 24728 45880 24734 45892
rect 25038 45880 25044 45892
rect 24728 45852 25044 45880
rect 24728 45840 24734 45852
rect 25038 45840 25044 45852
rect 25096 45840 25102 45892
rect 25148 45812 25176 45988
rect 25774 45948 25780 45960
rect 25735 45920 25780 45948
rect 25774 45908 25780 45920
rect 25832 45908 25838 45960
rect 25884 45948 25912 45988
rect 29914 45976 29920 45988
rect 29972 45976 29978 46028
rect 32030 46016 32036 46028
rect 31991 45988 32036 46016
rect 32030 45976 32036 45988
rect 32088 45976 32094 46028
rect 50614 46016 50620 46028
rect 33888 45988 36124 46016
rect 50575 45988 50620 46016
rect 28537 45951 28595 45957
rect 25884 45920 26234 45948
rect 25498 45840 25504 45892
rect 25556 45880 25562 45892
rect 26022 45883 26080 45889
rect 26022 45880 26034 45883
rect 25556 45852 26034 45880
rect 25556 45840 25562 45852
rect 26022 45849 26034 45852
rect 26068 45849 26080 45883
rect 26206 45880 26234 45920
rect 28537 45917 28549 45951
rect 28583 45948 28595 45951
rect 29822 45948 29828 45960
rect 28583 45920 29828 45948
rect 28583 45917 28595 45920
rect 28537 45911 28595 45917
rect 29822 45908 29828 45920
rect 29880 45908 29886 45960
rect 30184 45951 30242 45957
rect 30184 45917 30196 45951
rect 30230 45948 30242 45951
rect 30742 45948 30748 45960
rect 30230 45920 30748 45948
rect 30230 45917 30242 45920
rect 30184 45911 30242 45917
rect 30742 45908 30748 45920
rect 30800 45908 30806 45960
rect 33888 45948 33916 45988
rect 34054 45948 34060 45960
rect 30852 45920 33916 45948
rect 34015 45920 34060 45948
rect 28902 45880 28908 45892
rect 26206 45852 28908 45880
rect 26022 45843 26080 45849
rect 28902 45840 28908 45852
rect 28960 45840 28966 45892
rect 29362 45840 29368 45892
rect 29420 45880 29426 45892
rect 30852 45880 30880 45920
rect 34054 45908 34060 45920
rect 34112 45908 34118 45960
rect 34701 45951 34759 45957
rect 34701 45917 34713 45951
rect 34747 45948 34759 45951
rect 34790 45948 34796 45960
rect 34747 45920 34796 45948
rect 34747 45917 34759 45920
rect 34701 45911 34759 45917
rect 34790 45908 34796 45920
rect 34848 45908 34854 45960
rect 35526 45908 35532 45960
rect 35584 45948 35590 45960
rect 35805 45951 35863 45957
rect 35805 45948 35817 45951
rect 35584 45920 35817 45948
rect 35584 45908 35590 45920
rect 35805 45917 35817 45920
rect 35851 45917 35863 45951
rect 35805 45911 35863 45917
rect 29420 45852 30880 45880
rect 32300 45883 32358 45889
rect 29420 45840 29426 45852
rect 32300 45849 32312 45883
rect 32346 45880 32358 45883
rect 32346 45852 33916 45880
rect 32346 45849 32358 45852
rect 32300 45843 32358 45849
rect 23768 45784 25176 45812
rect 25590 45772 25596 45824
rect 25648 45812 25654 45824
rect 27157 45815 27215 45821
rect 27157 45812 27169 45815
rect 25648 45784 27169 45812
rect 25648 45772 25654 45784
rect 27157 45781 27169 45784
rect 27203 45781 27215 45815
rect 28350 45812 28356 45824
rect 28311 45784 28356 45812
rect 27157 45775 27215 45781
rect 28350 45772 28356 45784
rect 28408 45772 28414 45824
rect 30466 45772 30472 45824
rect 30524 45812 30530 45824
rect 31297 45815 31355 45821
rect 31297 45812 31309 45815
rect 30524 45784 31309 45812
rect 30524 45772 30530 45784
rect 31297 45781 31309 45784
rect 31343 45781 31355 45815
rect 31297 45775 31355 45781
rect 32674 45772 32680 45824
rect 32732 45812 32738 45824
rect 33888 45821 33916 45852
rect 34606 45840 34612 45892
rect 34664 45880 34670 45892
rect 35069 45883 35127 45889
rect 35069 45880 35081 45883
rect 34664 45852 35081 45880
rect 34664 45840 34670 45852
rect 35069 45849 35081 45852
rect 35115 45849 35127 45883
rect 35069 45843 35127 45849
rect 33413 45815 33471 45821
rect 33413 45812 33425 45815
rect 32732 45784 33425 45812
rect 32732 45772 32738 45784
rect 33413 45781 33425 45784
rect 33459 45781 33471 45815
rect 33413 45775 33471 45781
rect 33873 45815 33931 45821
rect 33873 45781 33885 45815
rect 33919 45781 33931 45815
rect 33873 45775 33931 45781
rect 35253 45815 35311 45821
rect 35253 45781 35265 45815
rect 35299 45812 35311 45815
rect 35618 45812 35624 45824
rect 35299 45784 35624 45812
rect 35299 45781 35311 45784
rect 35253 45775 35311 45781
rect 35618 45772 35624 45784
rect 35676 45772 35682 45824
rect 36096 45821 36124 45988
rect 50614 45976 50620 45988
rect 50672 45976 50678 46028
rect 40034 45948 40040 45960
rect 39995 45920 40040 45948
rect 40034 45908 40040 45920
rect 40092 45908 40098 45960
rect 40126 45908 40132 45960
rect 40184 45948 40190 45960
rect 40293 45951 40351 45957
rect 40293 45948 40305 45951
rect 40184 45920 40305 45948
rect 40184 45908 40190 45920
rect 40293 45917 40305 45920
rect 40339 45917 40351 45951
rect 42058 45948 42064 45960
rect 42019 45920 42064 45948
rect 40293 45911 40351 45917
rect 42058 45908 42064 45920
rect 42116 45908 42122 45960
rect 42150 45908 42156 45960
rect 42208 45948 42214 45960
rect 42317 45951 42375 45957
rect 42317 45948 42329 45951
rect 42208 45920 42329 45948
rect 42208 45908 42214 45920
rect 42317 45917 42329 45920
rect 42363 45917 42375 45951
rect 42317 45911 42375 45917
rect 45005 45951 45063 45957
rect 45005 45917 45017 45951
rect 45051 45917 45063 45951
rect 45005 45911 45063 45917
rect 45281 45951 45339 45957
rect 45281 45917 45293 45951
rect 45327 45948 45339 45951
rect 45741 45951 45799 45957
rect 45741 45948 45753 45951
rect 45327 45920 45753 45948
rect 45327 45917 45339 45920
rect 45281 45911 45339 45917
rect 45741 45917 45753 45920
rect 45787 45948 45799 45951
rect 46382 45948 46388 45960
rect 45787 45920 46388 45948
rect 45787 45917 45799 45920
rect 45741 45911 45799 45917
rect 36446 45840 36452 45892
rect 36504 45880 36510 45892
rect 36725 45883 36783 45889
rect 36725 45880 36737 45883
rect 36504 45852 36737 45880
rect 36504 45840 36510 45852
rect 36725 45849 36737 45852
rect 36771 45849 36783 45883
rect 45020 45880 45048 45911
rect 46382 45908 46388 45920
rect 46440 45908 46446 45960
rect 48038 45948 48044 45960
rect 47999 45920 48044 45948
rect 48038 45908 48044 45920
rect 48096 45908 48102 45960
rect 50801 45951 50859 45957
rect 50801 45917 50813 45951
rect 50847 45917 50859 45951
rect 50801 45911 50859 45917
rect 50985 45951 51043 45957
rect 50985 45917 50997 45951
rect 51031 45948 51043 45951
rect 51629 45951 51687 45957
rect 51629 45948 51641 45951
rect 51031 45920 51641 45948
rect 51031 45917 51043 45920
rect 50985 45911 51043 45917
rect 51629 45917 51641 45920
rect 51675 45917 51687 45951
rect 51629 45911 51687 45917
rect 45830 45880 45836 45892
rect 45020 45852 45836 45880
rect 36725 45843 36783 45849
rect 45830 45840 45836 45852
rect 45888 45840 45894 45892
rect 50816 45880 50844 45911
rect 66806 45908 66812 45960
rect 66864 45948 66870 45960
rect 67269 45951 67327 45957
rect 67269 45948 67281 45951
rect 66864 45920 67281 45948
rect 66864 45908 66870 45920
rect 67269 45917 67281 45920
rect 67315 45917 67327 45951
rect 67269 45911 67327 45917
rect 51718 45880 51724 45892
rect 50816 45852 51724 45880
rect 51718 45840 51724 45852
rect 51776 45840 51782 45892
rect 36081 45815 36139 45821
rect 36081 45781 36093 45815
rect 36127 45812 36139 45815
rect 37734 45812 37740 45824
rect 36127 45784 37740 45812
rect 36127 45781 36139 45784
rect 36081 45775 36139 45781
rect 37734 45772 37740 45784
rect 37792 45772 37798 45824
rect 51442 45812 51448 45824
rect 51403 45784 51448 45812
rect 51442 45772 51448 45784
rect 51500 45772 51506 45824
rect 1104 45722 68816 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 68816 45722
rect 1104 45648 68816 45670
rect 16574 45568 16580 45620
rect 16632 45608 16638 45620
rect 16853 45611 16911 45617
rect 16853 45608 16865 45611
rect 16632 45580 16865 45608
rect 16632 45568 16638 45580
rect 16853 45577 16865 45580
rect 16899 45577 16911 45611
rect 19242 45608 19248 45620
rect 16853 45571 16911 45577
rect 17696 45580 19248 45608
rect 12796 45543 12854 45549
rect 12796 45509 12808 45543
rect 12842 45540 12854 45543
rect 12986 45540 12992 45552
rect 12842 45512 12992 45540
rect 12842 45509 12854 45512
rect 12796 45503 12854 45509
rect 12986 45500 12992 45512
rect 13044 45500 13050 45552
rect 14820 45543 14878 45549
rect 14820 45509 14832 45543
rect 14866 45540 14878 45543
rect 15194 45540 15200 45552
rect 14866 45512 15200 45540
rect 14866 45509 14878 45512
rect 14820 45503 14878 45509
rect 15194 45500 15200 45512
rect 15252 45500 15258 45552
rect 1854 45472 1860 45484
rect 1815 45444 1860 45472
rect 1854 45432 1860 45444
rect 1912 45432 1918 45484
rect 14553 45475 14611 45481
rect 14553 45441 14565 45475
rect 14599 45472 14611 45475
rect 14642 45472 14648 45484
rect 14599 45444 14648 45472
rect 14599 45441 14611 45444
rect 14553 45435 14611 45441
rect 14642 45432 14648 45444
rect 14700 45432 14706 45484
rect 16853 45475 16911 45481
rect 16853 45441 16865 45475
rect 16899 45472 16911 45475
rect 16942 45472 16948 45484
rect 16899 45444 16948 45472
rect 16899 45441 16911 45444
rect 16853 45435 16911 45441
rect 16942 45432 16948 45444
rect 17000 45432 17006 45484
rect 17402 45432 17408 45484
rect 17460 45472 17466 45484
rect 17696 45481 17724 45580
rect 19242 45568 19248 45580
rect 19300 45568 19306 45620
rect 20622 45568 20628 45620
rect 20680 45608 20686 45620
rect 22278 45608 22284 45620
rect 20680 45580 22048 45608
rect 22239 45580 22284 45608
rect 20680 45568 20686 45580
rect 19337 45543 19395 45549
rect 19337 45509 19349 45543
rect 19383 45540 19395 45543
rect 21358 45540 21364 45552
rect 19383 45512 21364 45540
rect 19383 45509 19395 45512
rect 19337 45503 19395 45509
rect 21358 45500 21364 45512
rect 21416 45500 21422 45552
rect 21913 45543 21971 45549
rect 21913 45509 21925 45543
rect 21959 45509 21971 45543
rect 22020 45540 22048 45580
rect 22278 45568 22284 45580
rect 22336 45568 22342 45620
rect 24670 45608 24676 45620
rect 24631 45580 24676 45608
rect 24670 45568 24676 45580
rect 24728 45568 24734 45620
rect 24762 45568 24768 45620
rect 24820 45608 24826 45620
rect 29362 45608 29368 45620
rect 24820 45580 29368 45608
rect 24820 45568 24826 45580
rect 29362 45568 29368 45580
rect 29420 45568 29426 45620
rect 29822 45608 29828 45620
rect 29783 45580 29828 45608
rect 29822 45568 29828 45580
rect 29880 45568 29886 45620
rect 30745 45611 30803 45617
rect 30745 45577 30757 45611
rect 30791 45608 30803 45611
rect 30926 45608 30932 45620
rect 30791 45580 30932 45608
rect 30791 45577 30803 45580
rect 30745 45571 30803 45577
rect 30926 45568 30932 45580
rect 30984 45568 30990 45620
rect 42058 45568 42064 45620
rect 42116 45608 42122 45620
rect 42613 45611 42671 45617
rect 42613 45608 42625 45611
rect 42116 45580 42625 45608
rect 42116 45568 42122 45580
rect 42613 45577 42625 45580
rect 42659 45577 42671 45611
rect 42613 45571 42671 45577
rect 45373 45611 45431 45617
rect 45373 45577 45385 45611
rect 45419 45577 45431 45611
rect 45373 45571 45431 45577
rect 22113 45543 22171 45549
rect 22113 45540 22125 45543
rect 22020 45512 22125 45540
rect 21913 45503 21971 45509
rect 22113 45509 22125 45512
rect 22159 45509 22171 45543
rect 22113 45503 22171 45509
rect 23560 45543 23618 45549
rect 23560 45509 23572 45543
rect 23606 45540 23618 45543
rect 23658 45540 23664 45552
rect 23606 45512 23664 45540
rect 23606 45509 23618 45512
rect 23560 45503 23618 45509
rect 17497 45475 17555 45481
rect 17497 45472 17509 45475
rect 17460 45444 17509 45472
rect 17460 45432 17466 45444
rect 17497 45441 17509 45444
rect 17543 45441 17555 45475
rect 17497 45435 17555 45441
rect 17681 45475 17739 45481
rect 17681 45441 17693 45475
rect 17727 45441 17739 45475
rect 17681 45435 17739 45441
rect 18414 45432 18420 45484
rect 18472 45472 18478 45484
rect 20070 45481 20076 45484
rect 18472 45444 18517 45472
rect 18472 45432 18478 45444
rect 20064 45435 20076 45481
rect 20128 45472 20134 45484
rect 20128 45444 20164 45472
rect 20070 45432 20076 45435
rect 20128 45432 20134 45444
rect 21266 45432 21272 45484
rect 21324 45472 21330 45484
rect 21634 45472 21640 45484
rect 21324 45444 21640 45472
rect 21324 45432 21330 45444
rect 21634 45432 21640 45444
rect 21692 45472 21698 45484
rect 21928 45472 21956 45503
rect 23658 45500 23664 45512
rect 23716 45500 23722 45552
rect 24854 45500 24860 45552
rect 24912 45540 24918 45552
rect 25590 45540 25596 45552
rect 24912 45512 25596 45540
rect 24912 45500 24918 45512
rect 25590 45500 25596 45512
rect 25648 45500 25654 45552
rect 25682 45500 25688 45552
rect 25740 45540 25746 45552
rect 25793 45543 25851 45549
rect 25793 45540 25805 45543
rect 25740 45512 25805 45540
rect 25740 45500 25746 45512
rect 25793 45509 25805 45512
rect 25839 45509 25851 45543
rect 25793 45503 25851 45509
rect 27884 45543 27942 45549
rect 27884 45509 27896 45543
rect 27930 45540 27942 45543
rect 28350 45540 28356 45552
rect 27930 45512 28356 45540
rect 27930 45509 27942 45512
rect 27884 45503 27942 45509
rect 28350 45500 28356 45512
rect 28408 45500 28414 45552
rect 28810 45500 28816 45552
rect 28868 45540 28874 45552
rect 29457 45543 29515 45549
rect 29457 45540 29469 45543
rect 28868 45512 29469 45540
rect 28868 45500 28874 45512
rect 29457 45509 29469 45512
rect 29503 45509 29515 45543
rect 29457 45503 29515 45509
rect 29673 45543 29731 45549
rect 29673 45509 29685 45543
rect 29719 45540 29731 45543
rect 30377 45543 30435 45549
rect 29719 45512 30328 45540
rect 29719 45509 29731 45512
rect 29673 45503 29731 45509
rect 26970 45472 26976 45484
rect 21692 45444 21956 45472
rect 26931 45444 26976 45472
rect 21692 45432 21698 45444
rect 26970 45432 26976 45444
rect 27028 45432 27034 45484
rect 30300 45472 30328 45512
rect 30377 45509 30389 45543
rect 30423 45540 30435 45543
rect 30466 45540 30472 45552
rect 30423 45512 30472 45540
rect 30423 45509 30435 45512
rect 30377 45503 30435 45509
rect 30466 45500 30472 45512
rect 30524 45500 30530 45552
rect 30558 45500 30564 45552
rect 30616 45549 30622 45552
rect 30616 45543 30651 45549
rect 30639 45540 30651 45543
rect 32674 45540 32680 45552
rect 30639 45512 31754 45540
rect 32635 45512 32680 45540
rect 30639 45509 30651 45512
rect 30616 45503 30651 45509
rect 30616 45500 30622 45503
rect 30576 45472 30604 45500
rect 27448 45444 29592 45472
rect 30300 45444 30604 45472
rect 31726 45472 31754 45512
rect 32674 45500 32680 45512
rect 32732 45500 32738 45552
rect 32893 45543 32951 45549
rect 32893 45540 32905 45543
rect 32784 45512 32905 45540
rect 32784 45472 32812 45512
rect 32893 45509 32905 45512
rect 32939 45540 32951 45543
rect 34514 45540 34520 45552
rect 32939 45512 34520 45540
rect 32939 45509 32951 45512
rect 32893 45503 32951 45509
rect 34514 45500 34520 45512
rect 34572 45500 34578 45552
rect 34698 45500 34704 45552
rect 34756 45540 34762 45552
rect 37458 45540 37464 45552
rect 34756 45512 37320 45540
rect 34756 45500 34762 45512
rect 31726 45444 32812 45472
rect 34149 45475 34207 45481
rect 12526 45404 12532 45416
rect 12487 45376 12532 45404
rect 12526 45364 12532 45376
rect 12584 45364 12590 45416
rect 18534 45407 18592 45413
rect 18534 45404 18546 45407
rect 16546 45376 18546 45404
rect 16546 45336 16574 45376
rect 18534 45373 18546 45376
rect 18580 45373 18592 45407
rect 18534 45367 18592 45373
rect 18693 45407 18751 45413
rect 18693 45373 18705 45407
rect 18739 45404 18751 45407
rect 19058 45404 19064 45416
rect 18739 45376 19064 45404
rect 18739 45373 18751 45376
rect 18693 45367 18751 45373
rect 19058 45364 19064 45376
rect 19116 45364 19122 45416
rect 19426 45364 19432 45416
rect 19484 45404 19490 45416
rect 19797 45407 19855 45413
rect 19797 45404 19809 45407
rect 19484 45376 19809 45404
rect 19484 45364 19490 45376
rect 19797 45373 19809 45376
rect 19843 45373 19855 45407
rect 23290 45404 23296 45416
rect 23251 45376 23296 45404
rect 19797 45367 19855 45373
rect 23290 45364 23296 45376
rect 23348 45364 23354 45416
rect 25774 45364 25780 45416
rect 25832 45404 25838 45416
rect 27065 45407 27123 45413
rect 27065 45404 27077 45407
rect 25832 45376 27077 45404
rect 25832 45364 25838 45376
rect 27065 45373 27077 45376
rect 27111 45373 27123 45407
rect 27065 45367 27123 45373
rect 15488 45308 16574 45336
rect 18141 45339 18199 45345
rect 1946 45268 1952 45280
rect 1907 45240 1952 45268
rect 1946 45228 1952 45240
rect 2004 45228 2010 45280
rect 13170 45228 13176 45280
rect 13228 45268 13234 45280
rect 13909 45271 13967 45277
rect 13909 45268 13921 45271
rect 13228 45240 13921 45268
rect 13228 45228 13234 45240
rect 13909 45237 13921 45240
rect 13955 45268 13967 45271
rect 15488 45268 15516 45308
rect 18141 45305 18153 45339
rect 18187 45336 18199 45339
rect 18230 45336 18236 45348
rect 18187 45308 18236 45336
rect 18187 45305 18199 45308
rect 18141 45299 18199 45305
rect 18230 45296 18236 45308
rect 18288 45296 18294 45348
rect 27448 45336 27476 45444
rect 27614 45404 27620 45416
rect 27575 45376 27620 45404
rect 27614 45364 27620 45376
rect 27672 45364 27678 45416
rect 25792 45308 27476 45336
rect 15930 45268 15936 45280
rect 13955 45240 15516 45268
rect 15891 45240 15936 45268
rect 13955 45237 13967 45240
rect 13909 45231 13967 45237
rect 15930 45228 15936 45240
rect 15988 45268 15994 45280
rect 18414 45268 18420 45280
rect 15988 45240 18420 45268
rect 15988 45228 15994 45240
rect 18414 45228 18420 45240
rect 18472 45228 18478 45280
rect 20530 45228 20536 45280
rect 20588 45268 20594 45280
rect 25792 45277 25820 45308
rect 21177 45271 21235 45277
rect 21177 45268 21189 45271
rect 20588 45240 21189 45268
rect 20588 45228 20594 45240
rect 21177 45237 21189 45240
rect 21223 45237 21235 45271
rect 21177 45231 21235 45237
rect 22097 45271 22155 45277
rect 22097 45237 22109 45271
rect 22143 45268 22155 45271
rect 25777 45271 25835 45277
rect 25777 45268 25789 45271
rect 22143 45240 25789 45268
rect 22143 45237 22155 45240
rect 22097 45231 22155 45237
rect 25777 45237 25789 45240
rect 25823 45237 25835 45271
rect 25958 45268 25964 45280
rect 25919 45240 25964 45268
rect 25777 45231 25835 45237
rect 25958 45228 25964 45240
rect 26016 45228 26022 45280
rect 28810 45228 28816 45280
rect 28868 45268 28874 45280
rect 28997 45271 29055 45277
rect 28997 45268 29009 45271
rect 28868 45240 29009 45268
rect 28868 45228 28874 45240
rect 28997 45237 29009 45240
rect 29043 45237 29055 45271
rect 29564 45268 29592 45444
rect 34149 45441 34161 45475
rect 34195 45441 34207 45475
rect 35618 45472 35624 45484
rect 35579 45444 35624 45472
rect 34149 45435 34207 45441
rect 33045 45339 33103 45345
rect 33045 45305 33057 45339
rect 33091 45336 33103 45339
rect 34054 45336 34060 45348
rect 33091 45308 34060 45336
rect 33091 45305 33103 45308
rect 33045 45299 33103 45305
rect 34054 45296 34060 45308
rect 34112 45296 34118 45348
rect 34164 45336 34192 45435
rect 35618 45432 35624 45444
rect 35676 45432 35682 45484
rect 37292 45481 37320 45512
rect 37384 45512 37464 45540
rect 36449 45475 36507 45481
rect 36449 45441 36461 45475
rect 36495 45472 36507 45475
rect 37277 45475 37335 45481
rect 36495 45444 37228 45472
rect 36495 45441 36507 45444
rect 36449 45435 36507 45441
rect 34422 45404 34428 45416
rect 34383 45376 34428 45404
rect 34422 45364 34428 45376
rect 34480 45364 34486 45416
rect 34790 45364 34796 45416
rect 34848 45404 34854 45416
rect 36633 45407 36691 45413
rect 36633 45404 36645 45407
rect 34848 45376 36645 45404
rect 34848 45364 34854 45376
rect 36633 45373 36645 45376
rect 36679 45373 36691 45407
rect 36633 45367 36691 45373
rect 36725 45407 36783 45413
rect 36725 45373 36737 45407
rect 36771 45373 36783 45407
rect 37200 45404 37228 45444
rect 37277 45441 37289 45475
rect 37323 45441 37335 45475
rect 37277 45435 37335 45441
rect 37384 45404 37412 45512
rect 37458 45500 37464 45512
rect 37516 45500 37522 45552
rect 39384 45543 39442 45549
rect 39384 45509 39396 45543
rect 39430 45540 39442 45543
rect 39850 45540 39856 45552
rect 39430 45512 39856 45540
rect 39430 45509 39442 45512
rect 39384 45503 39442 45509
rect 39850 45500 39856 45512
rect 39908 45500 39914 45552
rect 43622 45500 43628 45552
rect 43680 45540 43686 45552
rect 45388 45540 45416 45571
rect 43680 45512 45416 45540
rect 50424 45543 50482 45549
rect 43680 45500 43686 45512
rect 50424 45509 50436 45543
rect 50470 45540 50482 45543
rect 51442 45540 51448 45552
rect 50470 45512 51448 45540
rect 50470 45509 50482 45512
rect 50424 45503 50482 45509
rect 51442 45500 51448 45512
rect 51500 45500 51506 45552
rect 37550 45481 37556 45484
rect 37544 45435 37556 45481
rect 37608 45472 37614 45484
rect 41141 45475 41199 45481
rect 37608 45444 37644 45472
rect 37550 45432 37556 45435
rect 37608 45432 37614 45444
rect 41141 45441 41153 45475
rect 41187 45472 41199 45475
rect 41414 45472 41420 45484
rect 41187 45444 41420 45472
rect 41187 45441 41199 45444
rect 41141 45435 41199 45441
rect 41414 45432 41420 45444
rect 41472 45472 41478 45484
rect 42429 45475 42487 45481
rect 42429 45472 42441 45475
rect 41472 45444 42441 45472
rect 41472 45432 41478 45444
rect 42429 45441 42441 45444
rect 42475 45441 42487 45475
rect 44910 45472 44916 45484
rect 44871 45444 44916 45472
rect 42429 45435 42487 45441
rect 44910 45432 44916 45444
rect 44968 45432 44974 45484
rect 45189 45475 45247 45481
rect 45189 45441 45201 45475
rect 45235 45472 45247 45475
rect 45646 45472 45652 45484
rect 45235 45444 45652 45472
rect 45235 45441 45247 45444
rect 45189 45435 45247 45441
rect 45646 45432 45652 45444
rect 45704 45432 45710 45484
rect 47765 45475 47823 45481
rect 47765 45441 47777 45475
rect 47811 45441 47823 45475
rect 47765 45435 47823 45441
rect 37200 45376 37412 45404
rect 39117 45407 39175 45413
rect 36725 45367 36783 45373
rect 39117 45373 39129 45407
rect 39163 45373 39175 45407
rect 39117 45367 39175 45373
rect 45097 45407 45155 45413
rect 45097 45373 45109 45407
rect 45143 45404 45155 45407
rect 45738 45404 45744 45416
rect 45143 45376 45744 45404
rect 45143 45373 45155 45376
rect 45097 45367 45155 45373
rect 35710 45336 35716 45348
rect 34164 45308 35716 45336
rect 35710 45296 35716 45308
rect 35768 45296 35774 45348
rect 29641 45271 29699 45277
rect 29641 45268 29653 45271
rect 29564 45240 29653 45268
rect 28997 45231 29055 45237
rect 29641 45237 29653 45240
rect 29687 45268 29699 45271
rect 30561 45271 30619 45277
rect 30561 45268 30573 45271
rect 29687 45240 30573 45268
rect 29687 45237 29699 45240
rect 29641 45231 29699 45237
rect 30561 45237 30573 45240
rect 30607 45268 30619 45271
rect 32858 45268 32864 45280
rect 30607 45240 32864 45268
rect 30607 45237 30619 45240
rect 30561 45231 30619 45237
rect 32858 45228 32864 45240
rect 32916 45228 32922 45280
rect 35434 45268 35440 45280
rect 35395 45240 35440 45268
rect 35434 45228 35440 45240
rect 35492 45228 35498 45280
rect 36262 45268 36268 45280
rect 36223 45240 36268 45268
rect 36262 45228 36268 45240
rect 36320 45228 36326 45280
rect 36740 45268 36768 45367
rect 37458 45268 37464 45280
rect 36740 45240 37464 45268
rect 37458 45228 37464 45240
rect 37516 45228 37522 45280
rect 38010 45228 38016 45280
rect 38068 45268 38074 45280
rect 38657 45271 38715 45277
rect 38657 45268 38669 45271
rect 38068 45240 38669 45268
rect 38068 45228 38074 45240
rect 38657 45237 38669 45240
rect 38703 45237 38715 45271
rect 39132 45268 39160 45367
rect 45738 45364 45744 45376
rect 45796 45364 45802 45416
rect 47780 45404 47808 45435
rect 47946 45432 47952 45484
rect 48004 45472 48010 45484
rect 48501 45475 48559 45481
rect 48501 45472 48513 45475
rect 48004 45444 48513 45472
rect 48004 45432 48010 45444
rect 48501 45441 48513 45444
rect 48547 45441 48559 45475
rect 48501 45435 48559 45441
rect 48038 45404 48044 45416
rect 47780 45376 48044 45404
rect 48038 45364 48044 45376
rect 48096 45404 48102 45416
rect 50154 45404 50160 45416
rect 48096 45376 48544 45404
rect 50115 45376 50160 45404
rect 48096 45364 48102 45376
rect 48516 45348 48544 45376
rect 50154 45364 50160 45376
rect 50212 45364 50218 45416
rect 40497 45339 40555 45345
rect 40497 45305 40509 45339
rect 40543 45336 40555 45339
rect 41506 45336 41512 45348
rect 40543 45308 41512 45336
rect 40543 45305 40555 45308
rect 40497 45299 40555 45305
rect 41506 45296 41512 45308
rect 41564 45296 41570 45348
rect 48498 45296 48504 45348
rect 48556 45296 48562 45348
rect 40957 45271 41015 45277
rect 40957 45268 40969 45271
rect 39132 45240 40969 45268
rect 38657 45231 38715 45237
rect 40957 45237 40969 45240
rect 41003 45237 41015 45271
rect 40957 45231 41015 45237
rect 45189 45271 45247 45277
rect 45189 45237 45201 45271
rect 45235 45268 45247 45271
rect 45554 45268 45560 45280
rect 45235 45240 45560 45268
rect 45235 45237 45247 45240
rect 45189 45231 45247 45237
rect 45554 45228 45560 45240
rect 45612 45228 45618 45280
rect 47578 45268 47584 45280
rect 47539 45240 47584 45268
rect 47578 45228 47584 45240
rect 47636 45228 47642 45280
rect 48314 45268 48320 45280
rect 48275 45240 48320 45268
rect 48314 45228 48320 45240
rect 48372 45228 48378 45280
rect 50798 45228 50804 45280
rect 50856 45268 50862 45280
rect 51537 45271 51595 45277
rect 51537 45268 51549 45271
rect 50856 45240 51549 45268
rect 50856 45228 50862 45240
rect 51537 45237 51549 45240
rect 51583 45237 51595 45271
rect 51537 45231 51595 45237
rect 66254 45228 66260 45280
rect 66312 45268 66318 45280
rect 67637 45271 67695 45277
rect 67637 45268 67649 45271
rect 66312 45240 67649 45268
rect 66312 45228 66318 45240
rect 67637 45237 67649 45240
rect 67683 45237 67695 45271
rect 67637 45231 67695 45237
rect 1104 45178 68816 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 65654 45178
rect 65706 45126 65718 45178
rect 65770 45126 65782 45178
rect 65834 45126 65846 45178
rect 65898 45126 65910 45178
rect 65962 45126 68816 45178
rect 1104 45104 68816 45126
rect 1946 45024 1952 45076
rect 2004 45064 2010 45076
rect 2004 45036 6914 45064
rect 2004 45024 2010 45036
rect 6886 44996 6914 45036
rect 12526 45024 12532 45076
rect 12584 45064 12590 45076
rect 12621 45067 12679 45073
rect 12621 45064 12633 45067
rect 12584 45036 12633 45064
rect 12584 45024 12590 45036
rect 12621 45033 12633 45036
rect 12667 45033 12679 45067
rect 13538 45064 13544 45076
rect 13499 45036 13544 45064
rect 12621 45027 12679 45033
rect 13538 45024 13544 45036
rect 13596 45024 13602 45076
rect 15470 45064 15476 45076
rect 15431 45036 15476 45064
rect 15470 45024 15476 45036
rect 15528 45024 15534 45076
rect 19426 45064 19432 45076
rect 19387 45036 19432 45064
rect 19426 45024 19432 45036
rect 19484 45024 19490 45076
rect 19981 45067 20039 45073
rect 19981 45033 19993 45067
rect 20027 45064 20039 45067
rect 20070 45064 20076 45076
rect 20027 45036 20076 45064
rect 20027 45033 20039 45036
rect 19981 45027 20039 45033
rect 20070 45024 20076 45036
rect 20128 45024 20134 45076
rect 21450 45064 21456 45076
rect 21411 45036 21456 45064
rect 21450 45024 21456 45036
rect 21508 45024 21514 45076
rect 25498 45024 25504 45076
rect 25556 45064 25562 45076
rect 25777 45067 25835 45073
rect 25777 45064 25789 45067
rect 25556 45036 25789 45064
rect 25556 45024 25562 45036
rect 25777 45033 25789 45036
rect 25823 45033 25835 45067
rect 27614 45064 27620 45076
rect 27575 45036 27620 45064
rect 25777 45027 25835 45033
rect 27614 45024 27620 45036
rect 27672 45024 27678 45076
rect 28902 45064 28908 45076
rect 28815 45036 28908 45064
rect 28902 45024 28908 45036
rect 28960 45064 28966 45076
rect 30650 45064 30656 45076
rect 28960 45036 30656 45064
rect 28960 45024 28966 45036
rect 30650 45024 30656 45036
rect 30708 45024 30714 45076
rect 37461 45067 37519 45073
rect 37461 45033 37473 45067
rect 37507 45064 37519 45067
rect 37550 45064 37556 45076
rect 37507 45036 37556 45064
rect 37507 45033 37519 45036
rect 37461 45027 37519 45033
rect 37550 45024 37556 45036
rect 37608 45024 37614 45076
rect 40034 45024 40040 45076
rect 40092 45064 40098 45076
rect 40129 45067 40187 45073
rect 40129 45064 40141 45067
rect 40092 45036 40141 45064
rect 40092 45024 40098 45036
rect 40129 45033 40141 45036
rect 40175 45033 40187 45067
rect 40129 45027 40187 45033
rect 45465 45067 45523 45073
rect 45465 45033 45477 45067
rect 45511 45064 45523 45067
rect 45554 45064 45560 45076
rect 45511 45036 45560 45064
rect 45511 45033 45523 45036
rect 45465 45027 45523 45033
rect 45554 45024 45560 45036
rect 45612 45064 45618 45076
rect 46658 45064 46664 45076
rect 45612 45036 46664 45064
rect 45612 45024 45618 45036
rect 46658 45024 46664 45036
rect 46716 45024 46722 45076
rect 50154 45064 50160 45076
rect 50115 45036 50160 45064
rect 50154 45024 50160 45036
rect 50212 45024 50218 45076
rect 19886 44996 19892 45008
rect 6886 44968 19892 44996
rect 19886 44956 19892 44968
rect 19944 44956 19950 45008
rect 30469 44999 30527 45005
rect 30469 44965 30481 44999
rect 30515 44996 30527 44999
rect 30558 44996 30564 45008
rect 30515 44968 30564 44996
rect 30515 44965 30527 44968
rect 30469 44959 30527 44965
rect 30558 44956 30564 44968
rect 30616 44956 30622 45008
rect 45649 44999 45707 45005
rect 45649 44965 45661 44999
rect 45695 44996 45707 44999
rect 46290 44996 46296 45008
rect 45695 44968 46296 44996
rect 45695 44965 45707 44968
rect 45649 44959 45707 44965
rect 46290 44956 46296 44968
rect 46348 44956 46354 45008
rect 13170 44928 13176 44940
rect 13131 44900 13176 44928
rect 13170 44888 13176 44900
rect 13228 44888 13234 44940
rect 15105 44931 15163 44937
rect 15105 44897 15117 44931
rect 15151 44928 15163 44931
rect 15930 44928 15936 44940
rect 15151 44900 15936 44928
rect 15151 44897 15163 44900
rect 15105 44891 15163 44897
rect 15930 44888 15936 44900
rect 15988 44888 15994 44940
rect 20806 44928 20812 44940
rect 19444 44900 20812 44928
rect 12618 44860 12624 44872
rect 12579 44832 12624 44860
rect 12618 44820 12624 44832
rect 12676 44820 12682 44872
rect 13354 44860 13360 44872
rect 13315 44832 13360 44860
rect 13354 44820 13360 44832
rect 13412 44820 13418 44872
rect 15286 44860 15292 44872
rect 15199 44832 15292 44860
rect 15286 44820 15292 44832
rect 15344 44860 15350 44872
rect 15562 44860 15568 44872
rect 15344 44832 15568 44860
rect 15344 44820 15350 44832
rect 15562 44820 15568 44832
rect 15620 44820 15626 44872
rect 19444 44869 19472 44900
rect 20806 44888 20812 44900
rect 20864 44888 20870 44940
rect 21082 44888 21088 44940
rect 21140 44928 21146 44940
rect 21140 44900 21956 44928
rect 21140 44888 21146 44900
rect 19429 44863 19487 44869
rect 19429 44829 19441 44863
rect 19475 44829 19487 44863
rect 19429 44823 19487 44829
rect 20165 44863 20223 44869
rect 20165 44829 20177 44863
rect 20211 44860 20223 44863
rect 20898 44860 20904 44872
rect 20211 44832 20904 44860
rect 20211 44829 20223 44832
rect 20165 44823 20223 44829
rect 20898 44820 20904 44832
rect 20956 44820 20962 44872
rect 21637 44863 21695 44869
rect 21637 44829 21649 44863
rect 21683 44860 21695 44863
rect 21818 44860 21824 44872
rect 21683 44832 21824 44860
rect 21683 44829 21695 44832
rect 21637 44823 21695 44829
rect 21818 44820 21824 44832
rect 21876 44820 21882 44872
rect 21928 44869 21956 44900
rect 26970 44888 26976 44940
rect 27028 44928 27034 44940
rect 30006 44928 30012 44940
rect 27028 44900 30012 44928
rect 27028 44888 27034 44900
rect 21913 44863 21971 44869
rect 21913 44829 21925 44863
rect 21959 44829 21971 44863
rect 21913 44823 21971 44829
rect 23017 44863 23075 44869
rect 23017 44829 23029 44863
rect 23063 44860 23075 44863
rect 23566 44860 23572 44872
rect 23063 44832 23572 44860
rect 23063 44829 23075 44832
rect 23017 44823 23075 44829
rect 23566 44820 23572 44832
rect 23624 44820 23630 44872
rect 25958 44860 25964 44872
rect 25919 44832 25964 44860
rect 25958 44820 25964 44832
rect 26016 44820 26022 44872
rect 27540 44869 27568 44900
rect 30006 44888 30012 44900
rect 30064 44888 30070 44940
rect 34698 44888 34704 44940
rect 34756 44928 34762 44940
rect 34885 44931 34943 44937
rect 34885 44928 34897 44931
rect 34756 44900 34897 44928
rect 34756 44888 34762 44900
rect 34885 44897 34897 44900
rect 34931 44897 34943 44931
rect 34885 44891 34943 44897
rect 38010 44888 38016 44940
rect 38068 44928 38074 44940
rect 38105 44931 38163 44937
rect 38105 44928 38117 44931
rect 38068 44900 38117 44928
rect 38068 44888 38074 44900
rect 38105 44897 38117 44900
rect 38151 44897 38163 44931
rect 44174 44928 44180 44940
rect 38105 44891 38163 44897
rect 42996 44900 44180 44928
rect 27525 44863 27583 44869
rect 27525 44829 27537 44863
rect 27571 44829 27583 44863
rect 27525 44823 27583 44829
rect 28350 44820 28356 44872
rect 28408 44860 28414 44872
rect 28721 44863 28779 44869
rect 28721 44860 28733 44863
rect 28408 44832 28733 44860
rect 28408 44820 28414 44832
rect 28721 44829 28733 44832
rect 28767 44829 28779 44863
rect 31110 44860 31116 44872
rect 31071 44832 31116 44860
rect 28721 44823 28779 44829
rect 31110 44820 31116 44832
rect 31168 44820 31174 44872
rect 32490 44860 32496 44872
rect 32451 44832 32496 44860
rect 32490 44820 32496 44832
rect 32548 44820 32554 44872
rect 35152 44863 35210 44869
rect 35152 44829 35164 44863
rect 35198 44860 35210 44863
rect 35434 44860 35440 44872
rect 35198 44832 35440 44860
rect 35198 44829 35210 44832
rect 35152 44823 35210 44829
rect 35434 44820 35440 44832
rect 35492 44820 35498 44872
rect 37645 44863 37703 44869
rect 37645 44829 37657 44863
rect 37691 44829 37703 44863
rect 37645 44823 37703 44829
rect 38289 44863 38347 44869
rect 38289 44829 38301 44863
rect 38335 44860 38347 44863
rect 40129 44863 40187 44869
rect 38335 44832 39896 44860
rect 38335 44829 38347 44832
rect 38289 44823 38347 44829
rect 20714 44752 20720 44804
rect 20772 44792 20778 44804
rect 23109 44795 23167 44801
rect 23109 44792 23121 44795
rect 20772 44764 23121 44792
rect 20772 44752 20778 44764
rect 23109 44761 23121 44764
rect 23155 44761 23167 44795
rect 23109 44755 23167 44761
rect 30006 44752 30012 44804
rect 30064 44792 30070 44804
rect 30282 44792 30288 44804
rect 30064 44764 30288 44792
rect 30064 44752 30070 44764
rect 30282 44752 30288 44764
rect 30340 44752 30346 44804
rect 37660 44792 37688 44823
rect 38473 44795 38531 44801
rect 38473 44792 38485 44795
rect 37660 44764 38485 44792
rect 38473 44761 38485 44764
rect 38519 44761 38531 44795
rect 39868 44792 39896 44832
rect 40129 44829 40141 44863
rect 40175 44860 40187 44863
rect 41414 44860 41420 44872
rect 40175 44832 41420 44860
rect 40175 44829 40187 44832
rect 40129 44823 40187 44829
rect 41414 44820 41420 44832
rect 41472 44820 41478 44872
rect 41690 44860 41696 44872
rect 41651 44832 41696 44860
rect 41690 44820 41696 44832
rect 41748 44820 41754 44872
rect 41782 44820 41788 44872
rect 41840 44860 41846 44872
rect 41949 44863 42007 44869
rect 41949 44860 41961 44863
rect 41840 44832 41961 44860
rect 41840 44820 41846 44832
rect 41949 44829 41961 44832
rect 41995 44829 42007 44863
rect 41949 44823 42007 44829
rect 42996 44792 43024 44900
rect 44174 44888 44180 44900
rect 44232 44888 44238 44940
rect 45373 44931 45431 44937
rect 45373 44897 45385 44931
rect 45419 44928 45431 44931
rect 45738 44928 45744 44940
rect 45419 44900 45744 44928
rect 45419 44897 45431 44900
rect 45373 44891 45431 44897
rect 45738 44888 45744 44900
rect 45796 44888 45802 44940
rect 47578 44928 47584 44940
rect 47539 44900 47584 44928
rect 47578 44888 47584 44900
rect 47636 44888 47642 44940
rect 66254 44928 66260 44940
rect 66215 44900 66260 44928
rect 66254 44888 66260 44900
rect 66312 44888 66318 44940
rect 68094 44928 68100 44940
rect 68055 44900 68100 44928
rect 68094 44888 68100 44900
rect 68152 44888 68158 44940
rect 43993 44863 44051 44869
rect 43993 44829 44005 44863
rect 44039 44860 44051 44863
rect 44358 44860 44364 44872
rect 44039 44832 44364 44860
rect 44039 44829 44051 44832
rect 43993 44823 44051 44829
rect 44358 44820 44364 44832
rect 44416 44820 44422 44872
rect 45465 44863 45523 44869
rect 45465 44829 45477 44863
rect 45511 44860 45523 44863
rect 45646 44860 45652 44872
rect 45511 44832 45652 44860
rect 45511 44829 45523 44832
rect 45465 44823 45523 44829
rect 45646 44820 45652 44832
rect 45704 44860 45710 44872
rect 46198 44860 46204 44872
rect 45704 44832 46204 44860
rect 45704 44820 45710 44832
rect 46198 44820 46204 44832
rect 46256 44820 46262 44872
rect 46293 44863 46351 44869
rect 46293 44829 46305 44863
rect 46339 44860 46351 44863
rect 47848 44863 47906 44869
rect 46339 44832 47808 44860
rect 46339 44829 46351 44832
rect 46293 44823 46351 44829
rect 43530 44792 43536 44804
rect 39868 44764 43024 44792
rect 43088 44764 43536 44792
rect 38473 44755 38531 44761
rect 21821 44727 21879 44733
rect 21821 44693 21833 44727
rect 21867 44724 21879 44727
rect 21910 44724 21916 44736
rect 21867 44696 21916 44724
rect 21867 44693 21879 44696
rect 21821 44687 21879 44693
rect 21910 44684 21916 44696
rect 21968 44684 21974 44736
rect 30926 44684 30932 44736
rect 30984 44724 30990 44736
rect 31113 44727 31171 44733
rect 31113 44724 31125 44727
rect 30984 44696 31125 44724
rect 30984 44684 30990 44696
rect 31113 44693 31125 44696
rect 31159 44693 31171 44727
rect 31113 44687 31171 44693
rect 32585 44727 32643 44733
rect 32585 44693 32597 44727
rect 32631 44724 32643 44727
rect 34330 44724 34336 44736
rect 32631 44696 34336 44724
rect 32631 44693 32643 44696
rect 32585 44687 32643 44693
rect 34330 44684 34336 44696
rect 34388 44684 34394 44736
rect 36170 44684 36176 44736
rect 36228 44724 36234 44736
rect 43088 44733 43116 44764
rect 43530 44752 43536 44764
rect 43588 44792 43594 44804
rect 45005 44795 45063 44801
rect 45005 44792 45017 44795
rect 43588 44764 45017 44792
rect 43588 44752 43594 44764
rect 45005 44761 45017 44764
rect 45051 44761 45063 44795
rect 47780 44792 47808 44832
rect 47848 44829 47860 44863
rect 47894 44860 47906 44863
rect 48314 44860 48320 44872
rect 47894 44832 48320 44860
rect 47894 44829 47906 44832
rect 47848 44823 47906 44829
rect 48314 44820 48320 44832
rect 48372 44820 48378 44872
rect 50341 44863 50399 44869
rect 50341 44829 50353 44863
rect 50387 44860 50399 44863
rect 51350 44860 51356 44872
rect 50387 44832 51356 44860
rect 50387 44829 50399 44832
rect 50341 44823 50399 44829
rect 51350 44820 51356 44832
rect 51408 44820 51414 44872
rect 48406 44792 48412 44804
rect 47780 44764 48412 44792
rect 45005 44755 45063 44761
rect 48406 44752 48412 44764
rect 48464 44752 48470 44804
rect 66438 44792 66444 44804
rect 66399 44764 66444 44792
rect 66438 44752 66444 44764
rect 66496 44752 66502 44804
rect 36265 44727 36323 44733
rect 36265 44724 36277 44727
rect 36228 44696 36277 44724
rect 36228 44684 36234 44696
rect 36265 44693 36277 44696
rect 36311 44693 36323 44727
rect 36265 44687 36323 44693
rect 43073 44727 43131 44733
rect 43073 44693 43085 44727
rect 43119 44693 43131 44727
rect 43806 44724 43812 44736
rect 43767 44696 43812 44724
rect 43073 44687 43131 44693
rect 43806 44684 43812 44696
rect 43864 44684 43870 44736
rect 44174 44684 44180 44736
rect 44232 44724 44238 44736
rect 46523 44727 46581 44733
rect 46523 44724 46535 44727
rect 44232 44696 46535 44724
rect 44232 44684 44238 44696
rect 46523 44693 46535 44696
rect 46569 44693 46581 44727
rect 46523 44687 46581 44693
rect 46658 44684 46664 44736
rect 46716 44724 46722 44736
rect 47670 44724 47676 44736
rect 46716 44696 47676 44724
rect 46716 44684 46722 44696
rect 47670 44684 47676 44696
rect 47728 44724 47734 44736
rect 48961 44727 49019 44733
rect 48961 44724 48973 44727
rect 47728 44696 48973 44724
rect 47728 44684 47734 44696
rect 48961 44693 48973 44696
rect 49007 44693 49019 44727
rect 48961 44687 49019 44693
rect 1104 44634 68816 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 68816 44634
rect 1104 44560 68816 44582
rect 14550 44480 14556 44532
rect 14608 44520 14614 44532
rect 14645 44523 14703 44529
rect 14645 44520 14657 44523
rect 14608 44492 14657 44520
rect 14608 44480 14614 44492
rect 14645 44489 14657 44492
rect 14691 44489 14703 44523
rect 20530 44520 20536 44532
rect 14645 44483 14703 44489
rect 18156 44492 20536 44520
rect 12618 44384 12624 44396
rect 12579 44356 12624 44384
rect 12618 44344 12624 44356
rect 12676 44344 12682 44396
rect 14461 44387 14519 44393
rect 14461 44353 14473 44387
rect 14507 44384 14519 44387
rect 14734 44384 14740 44396
rect 14507 44356 14740 44384
rect 14507 44353 14519 44356
rect 14461 44347 14519 44353
rect 14734 44344 14740 44356
rect 14792 44344 14798 44396
rect 15378 44384 15384 44396
rect 15339 44356 15384 44384
rect 15378 44344 15384 44356
rect 15436 44344 15442 44396
rect 16853 44387 16911 44393
rect 16853 44353 16865 44387
rect 16899 44384 16911 44387
rect 17034 44384 17040 44396
rect 16899 44356 17040 44384
rect 16899 44353 16911 44356
rect 16853 44347 16911 44353
rect 17034 44344 17040 44356
rect 17092 44344 17098 44396
rect 18156 44393 18184 44492
rect 20530 44480 20536 44492
rect 20588 44480 20594 44532
rect 23290 44480 23296 44532
rect 23348 44520 23354 44532
rect 23385 44523 23443 44529
rect 23385 44520 23397 44523
rect 23348 44492 23397 44520
rect 23348 44480 23354 44492
rect 23385 44489 23397 44492
rect 23431 44489 23443 44523
rect 23385 44483 23443 44489
rect 29914 44480 29920 44532
rect 29972 44520 29978 44532
rect 30945 44523 31003 44529
rect 30945 44520 30957 44523
rect 29972 44492 30957 44520
rect 29972 44480 29978 44492
rect 30945 44489 30957 44492
rect 30991 44489 31003 44523
rect 30945 44483 31003 44489
rect 31113 44523 31171 44529
rect 31113 44489 31125 44523
rect 31159 44489 31171 44523
rect 31113 44483 31171 44489
rect 21910 44412 21916 44464
rect 21968 44452 21974 44464
rect 22741 44455 22799 44461
rect 22741 44452 22753 44455
rect 21968 44424 22753 44452
rect 21968 44412 21974 44424
rect 22741 44421 22753 44424
rect 22787 44421 22799 44455
rect 24026 44452 24032 44464
rect 22741 44415 22799 44421
rect 22848 44424 24032 44452
rect 18141 44387 18199 44393
rect 18141 44353 18153 44387
rect 18187 44353 18199 44387
rect 18141 44347 18199 44353
rect 21818 44344 21824 44396
rect 21876 44384 21882 44396
rect 22848 44393 22876 44424
rect 24026 44412 24032 44424
rect 24084 44412 24090 44464
rect 30742 44452 30748 44464
rect 30703 44424 30748 44452
rect 30742 44412 30748 44424
rect 30800 44412 30806 44464
rect 22557 44387 22615 44393
rect 22557 44384 22569 44387
rect 21876 44356 22569 44384
rect 21876 44344 21882 44356
rect 22557 44353 22569 44356
rect 22603 44353 22615 44387
rect 22557 44347 22615 44353
rect 22833 44387 22891 44393
rect 22833 44353 22845 44387
rect 22879 44353 22891 44387
rect 22833 44347 22891 44353
rect 23293 44387 23351 44393
rect 23293 44353 23305 44387
rect 23339 44384 23351 44387
rect 23566 44384 23572 44396
rect 23339 44356 23572 44384
rect 23339 44353 23351 44356
rect 23293 44347 23351 44353
rect 23566 44344 23572 44356
rect 23624 44384 23630 44396
rect 25222 44384 25228 44396
rect 23624 44356 24072 44384
rect 25183 44356 25228 44384
rect 23624 44344 23630 44356
rect 24044 44328 24072 44356
rect 25222 44344 25228 44356
rect 25280 44344 25286 44396
rect 27157 44387 27215 44393
rect 27157 44353 27169 44387
rect 27203 44384 27215 44387
rect 28902 44384 28908 44396
rect 27203 44356 28908 44384
rect 27203 44353 27215 44356
rect 27157 44347 27215 44353
rect 28902 44344 28908 44356
rect 28960 44344 28966 44396
rect 30101 44387 30159 44393
rect 30101 44353 30113 44387
rect 30147 44353 30159 44387
rect 31128 44384 31156 44483
rect 34606 44480 34612 44532
rect 34664 44480 34670 44532
rect 34698 44480 34704 44532
rect 34756 44520 34762 44532
rect 34793 44523 34851 44529
rect 34793 44520 34805 44523
rect 34756 44492 34805 44520
rect 34756 44480 34762 44492
rect 34793 44489 34805 44492
rect 34839 44489 34851 44523
rect 34793 44483 34851 44489
rect 32309 44387 32367 44393
rect 32309 44384 32321 44387
rect 31128 44356 32321 44384
rect 30101 44347 30159 44353
rect 32309 44353 32321 44356
rect 32355 44353 32367 44387
rect 32309 44347 32367 44353
rect 33965 44387 34023 44393
rect 33965 44353 33977 44387
rect 34011 44384 34023 44387
rect 34146 44384 34152 44396
rect 34011 44356 34152 44384
rect 34011 44353 34023 44356
rect 33965 44347 34023 44353
rect 17954 44316 17960 44328
rect 17915 44288 17960 44316
rect 17954 44276 17960 44288
rect 18012 44276 18018 44328
rect 18877 44319 18935 44325
rect 18877 44316 18889 44319
rect 18248 44288 18889 44316
rect 16758 44208 16764 44260
rect 16816 44248 16822 44260
rect 18248 44248 18276 44288
rect 18877 44285 18889 44288
rect 18923 44285 18935 44319
rect 18877 44279 18935 44285
rect 18966 44276 18972 44328
rect 19024 44325 19030 44328
rect 19024 44319 19052 44325
rect 19040 44285 19052 44319
rect 19024 44279 19052 44285
rect 19024 44276 19030 44279
rect 19150 44276 19156 44328
rect 19208 44316 19214 44328
rect 19208 44288 19253 44316
rect 19208 44276 19214 44288
rect 24026 44276 24032 44328
rect 24084 44276 24090 44328
rect 30116 44316 30144 44347
rect 34146 44344 34152 44356
rect 34204 44344 34210 44396
rect 34624 44328 34652 44480
rect 34808 44452 34836 44483
rect 41690 44480 41696 44532
rect 41748 44520 41754 44532
rect 41785 44523 41843 44529
rect 41785 44520 41797 44523
rect 41748 44492 41797 44520
rect 41748 44480 41754 44492
rect 41785 44489 41797 44492
rect 41831 44489 41843 44523
rect 41785 44483 41843 44489
rect 44545 44523 44603 44529
rect 44545 44489 44557 44523
rect 44591 44520 44603 44523
rect 44910 44520 44916 44532
rect 44591 44492 44916 44520
rect 44591 44489 44603 44492
rect 44545 44483 44603 44489
rect 44910 44480 44916 44492
rect 44968 44480 44974 44532
rect 45830 44520 45836 44532
rect 45791 44492 45836 44520
rect 45830 44480 45836 44492
rect 45888 44480 45894 44532
rect 47946 44520 47952 44532
rect 47907 44492 47952 44520
rect 47946 44480 47952 44492
rect 48004 44480 48010 44532
rect 49421 44523 49479 44529
rect 49421 44489 49433 44523
rect 49467 44520 49479 44523
rect 51350 44520 51356 44532
rect 49467 44492 51356 44520
rect 49467 44489 49479 44492
rect 49421 44483 49479 44489
rect 51350 44480 51356 44492
rect 51408 44480 51414 44532
rect 66438 44480 66444 44532
rect 66496 44520 66502 44532
rect 67545 44523 67603 44529
rect 67545 44520 67557 44523
rect 66496 44492 67557 44520
rect 66496 44480 66502 44492
rect 67545 44489 67557 44492
rect 67591 44489 67603 44523
rect 67545 44483 67603 44489
rect 35612 44455 35670 44461
rect 34808 44424 35388 44452
rect 34701 44387 34759 44393
rect 34701 44353 34713 44387
rect 34747 44384 34759 44387
rect 34790 44384 34796 44396
rect 34747 44356 34796 44384
rect 34747 44353 34759 44356
rect 34701 44347 34759 44353
rect 34790 44344 34796 44356
rect 34848 44344 34854 44396
rect 35360 44393 35388 44424
rect 35612 44421 35624 44455
rect 35658 44452 35670 44455
rect 36262 44452 36268 44464
rect 35658 44424 36268 44452
rect 35658 44421 35670 44424
rect 35612 44415 35670 44421
rect 36262 44412 36268 44424
rect 36320 44412 36326 44464
rect 41046 44412 41052 44464
rect 41104 44452 41110 44464
rect 41104 44424 60734 44452
rect 41104 44412 41110 44424
rect 35345 44387 35403 44393
rect 35345 44353 35357 44387
rect 35391 44353 35403 44387
rect 35345 44347 35403 44353
rect 41414 44344 41420 44396
rect 41472 44384 41478 44396
rect 41601 44387 41659 44393
rect 41601 44384 41613 44387
rect 41472 44356 41613 44384
rect 41472 44344 41478 44356
rect 41601 44353 41613 44356
rect 41647 44353 41659 44387
rect 41601 44347 41659 44353
rect 42429 44387 42487 44393
rect 42429 44353 42441 44387
rect 42475 44384 42487 44387
rect 42518 44384 42524 44396
rect 42475 44356 42524 44384
rect 42475 44353 42487 44356
rect 42429 44347 42487 44353
rect 34514 44316 34520 44328
rect 30116 44288 34520 44316
rect 34514 44276 34520 44288
rect 34572 44276 34578 44328
rect 34606 44276 34612 44328
rect 34664 44276 34670 44328
rect 16816 44220 18276 44248
rect 16816 44208 16822 44220
rect 18322 44208 18328 44260
rect 18380 44248 18386 44260
rect 18601 44251 18659 44257
rect 18601 44248 18613 44251
rect 18380 44220 18613 44248
rect 18380 44208 18386 44220
rect 18601 44217 18613 44220
rect 18647 44217 18659 44251
rect 41616 44248 41644 44347
rect 42518 44344 42524 44356
rect 42576 44344 42582 44396
rect 43432 44387 43490 44393
rect 43432 44353 43444 44387
rect 43478 44384 43490 44387
rect 43806 44384 43812 44396
rect 43478 44356 43812 44384
rect 43478 44353 43490 44356
rect 43432 44347 43490 44353
rect 43806 44344 43812 44356
rect 43864 44344 43870 44396
rect 45465 44387 45523 44393
rect 45465 44353 45477 44387
rect 45511 44384 45523 44387
rect 45738 44384 45744 44396
rect 45511 44356 45744 44384
rect 45511 44353 45523 44356
rect 45465 44347 45523 44353
rect 45738 44344 45744 44356
rect 45796 44344 45802 44396
rect 46293 44387 46351 44393
rect 46293 44353 46305 44387
rect 46339 44353 46351 44387
rect 47670 44384 47676 44396
rect 47631 44356 47676 44384
rect 46293 44347 46351 44353
rect 43162 44316 43168 44328
rect 43123 44288 43168 44316
rect 43162 44276 43168 44288
rect 43220 44276 43226 44328
rect 45557 44319 45615 44325
rect 45557 44285 45569 44319
rect 45603 44316 45615 44319
rect 46198 44316 46204 44328
rect 45603 44288 46204 44316
rect 45603 44285 45615 44288
rect 45557 44279 45615 44285
rect 46198 44276 46204 44288
rect 46256 44276 46262 44328
rect 46308 44316 46336 44347
rect 47670 44344 47676 44356
rect 47728 44344 47734 44396
rect 47762 44344 47768 44396
rect 47820 44384 47826 44396
rect 48498 44384 48504 44396
rect 47820 44356 47865 44384
rect 48459 44356 48504 44384
rect 47820 44344 47826 44356
rect 48498 44344 48504 44356
rect 48556 44344 48562 44396
rect 48682 44344 48688 44396
rect 48740 44384 48746 44396
rect 49237 44387 49295 44393
rect 49237 44384 49249 44387
rect 48740 44356 49249 44384
rect 48740 44344 48746 44356
rect 49237 44353 49249 44356
rect 49283 44353 49295 44387
rect 60706 44384 60734 44424
rect 66622 44384 66628 44396
rect 60706 44356 66628 44384
rect 49237 44347 49295 44353
rect 66622 44344 66628 44356
rect 66680 44384 66686 44396
rect 67453 44387 67511 44393
rect 67453 44384 67465 44387
rect 66680 44356 67465 44384
rect 66680 44344 66686 44356
rect 67453 44353 67465 44356
rect 67499 44353 67511 44387
rect 67453 44347 67511 44353
rect 48516 44316 48544 44344
rect 46308 44288 48544 44316
rect 42426 44248 42432 44260
rect 41616 44220 42432 44248
rect 18601 44211 18659 44217
rect 42426 44208 42432 44220
rect 42484 44248 42490 44260
rect 42613 44251 42671 44257
rect 42613 44248 42625 44251
rect 42484 44220 42625 44248
rect 42484 44208 42490 44220
rect 42613 44217 42625 44220
rect 42659 44217 42671 44251
rect 42613 44211 42671 44217
rect 45646 44208 45652 44260
rect 45704 44248 45710 44260
rect 46385 44251 46443 44257
rect 46385 44248 46397 44251
rect 45704 44220 46397 44248
rect 45704 44208 45710 44220
rect 46385 44217 46397 44220
rect 46431 44217 46443 44251
rect 46385 44211 46443 44217
rect 12618 44180 12624 44192
rect 12579 44152 12624 44180
rect 12618 44140 12624 44152
rect 12676 44140 12682 44192
rect 15194 44180 15200 44192
rect 15155 44152 15200 44180
rect 15194 44140 15200 44152
rect 15252 44140 15258 44192
rect 16669 44183 16727 44189
rect 16669 44149 16681 44183
rect 16715 44180 16727 44183
rect 16850 44180 16856 44192
rect 16715 44152 16856 44180
rect 16715 44149 16727 44152
rect 16669 44143 16727 44149
rect 16850 44140 16856 44152
rect 16908 44140 16914 44192
rect 19797 44183 19855 44189
rect 19797 44149 19809 44183
rect 19843 44180 19855 44183
rect 20990 44180 20996 44192
rect 19843 44152 20996 44180
rect 19843 44149 19855 44152
rect 19797 44143 19855 44149
rect 20990 44140 20996 44152
rect 21048 44140 21054 44192
rect 22002 44140 22008 44192
rect 22060 44180 22066 44192
rect 22373 44183 22431 44189
rect 22373 44180 22385 44183
rect 22060 44152 22385 44180
rect 22060 44140 22066 44152
rect 22373 44149 22385 44152
rect 22419 44149 22431 44183
rect 25038 44180 25044 44192
rect 24999 44152 25044 44180
rect 22373 44143 22431 44149
rect 25038 44140 25044 44152
rect 25096 44140 25102 44192
rect 26973 44183 27031 44189
rect 26973 44149 26985 44183
rect 27019 44180 27031 44183
rect 27246 44180 27252 44192
rect 27019 44152 27252 44180
rect 27019 44149 27031 44152
rect 26973 44143 27031 44149
rect 27246 44140 27252 44152
rect 27304 44140 27310 44192
rect 28350 44140 28356 44192
rect 28408 44180 28414 44192
rect 30193 44183 30251 44189
rect 30193 44180 30205 44183
rect 28408 44152 30205 44180
rect 28408 44140 28414 44152
rect 30193 44149 30205 44152
rect 30239 44180 30251 44183
rect 30558 44180 30564 44192
rect 30239 44152 30564 44180
rect 30239 44149 30251 44152
rect 30193 44143 30251 44149
rect 30558 44140 30564 44152
rect 30616 44140 30622 44192
rect 30929 44183 30987 44189
rect 30929 44149 30941 44183
rect 30975 44180 30987 44183
rect 31202 44180 31208 44192
rect 30975 44152 31208 44180
rect 30975 44149 30987 44152
rect 30929 44143 30987 44149
rect 31202 44140 31208 44152
rect 31260 44140 31266 44192
rect 32122 44180 32128 44192
rect 32083 44152 32128 44180
rect 32122 44140 32128 44152
rect 32180 44140 32186 44192
rect 33778 44180 33784 44192
rect 33739 44152 33784 44180
rect 33778 44140 33784 44152
rect 33836 44140 33842 44192
rect 36262 44140 36268 44192
rect 36320 44180 36326 44192
rect 36725 44183 36783 44189
rect 36725 44180 36737 44183
rect 36320 44152 36737 44180
rect 36320 44140 36326 44152
rect 36725 44149 36737 44152
rect 36771 44149 36783 44183
rect 36725 44143 36783 44149
rect 45465 44183 45523 44189
rect 45465 44149 45477 44183
rect 45511 44180 45523 44183
rect 45554 44180 45560 44192
rect 45511 44152 45560 44180
rect 45511 44149 45523 44152
rect 45465 44143 45523 44149
rect 45554 44140 45560 44152
rect 45612 44140 45618 44192
rect 48590 44180 48596 44192
rect 48551 44152 48596 44180
rect 48590 44140 48596 44152
rect 48648 44140 48654 44192
rect 1104 44090 68816 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 65654 44090
rect 65706 44038 65718 44090
rect 65770 44038 65782 44090
rect 65834 44038 65846 44090
rect 65898 44038 65910 44090
rect 65962 44038 68816 44090
rect 1104 44016 68816 44038
rect 1949 43979 2007 43985
rect 1949 43945 1961 43979
rect 1995 43976 2007 43979
rect 20530 43976 20536 43988
rect 1995 43948 20536 43976
rect 1995 43945 2007 43948
rect 1949 43939 2007 43945
rect 20530 43936 20536 43948
rect 20588 43936 20594 43988
rect 28994 43976 29000 43988
rect 20916 43948 29000 43976
rect 16025 43911 16083 43917
rect 16025 43877 16037 43911
rect 16071 43908 16083 43911
rect 16574 43908 16580 43920
rect 16071 43880 16580 43908
rect 16071 43877 16083 43880
rect 16025 43871 16083 43877
rect 16574 43868 16580 43880
rect 16632 43908 16638 43920
rect 16758 43908 16764 43920
rect 16632 43880 16764 43908
rect 16632 43868 16638 43880
rect 16758 43868 16764 43880
rect 16816 43868 16822 43920
rect 18322 43868 18328 43920
rect 18380 43908 18386 43920
rect 19058 43908 19064 43920
rect 18380 43880 19064 43908
rect 18380 43868 18386 43880
rect 19058 43868 19064 43880
rect 19116 43908 19122 43920
rect 20349 43911 20407 43917
rect 20349 43908 20361 43911
rect 19116 43880 20361 43908
rect 19116 43868 19122 43880
rect 20349 43877 20361 43880
rect 20395 43877 20407 43911
rect 20349 43871 20407 43877
rect 13265 43775 13323 43781
rect 13265 43741 13277 43775
rect 13311 43741 13323 43775
rect 13265 43735 13323 43741
rect 1854 43704 1860 43716
rect 1815 43676 1860 43704
rect 1854 43664 1860 43676
rect 1912 43664 1918 43716
rect 13280 43704 13308 43735
rect 13354 43732 13360 43784
rect 13412 43772 13418 43784
rect 14642 43772 14648 43784
rect 13412 43744 14228 43772
rect 14603 43744 14648 43772
rect 13412 43732 13418 43744
rect 14090 43704 14096 43716
rect 13280 43676 14096 43704
rect 14090 43664 14096 43676
rect 14148 43664 14154 43716
rect 14200 43704 14228 43744
rect 14642 43732 14648 43744
rect 14700 43732 14706 43784
rect 14912 43775 14970 43781
rect 14912 43741 14924 43775
rect 14958 43772 14970 43775
rect 15194 43772 15200 43784
rect 14958 43744 15200 43772
rect 14958 43741 14970 43744
rect 14912 43735 14970 43741
rect 15194 43732 15200 43744
rect 15252 43732 15258 43784
rect 16761 43775 16819 43781
rect 16761 43741 16773 43775
rect 16807 43741 16819 43775
rect 16761 43735 16819 43741
rect 15746 43704 15752 43716
rect 14200 43676 15752 43704
rect 15746 43664 15752 43676
rect 15804 43664 15810 43716
rect 16776 43704 16804 43735
rect 16850 43732 16856 43784
rect 16908 43772 16914 43784
rect 17017 43775 17075 43781
rect 17017 43772 17029 43775
rect 16908 43744 17029 43772
rect 16908 43732 16914 43744
rect 17017 43741 17029 43744
rect 17063 43741 17075 43775
rect 17017 43735 17075 43741
rect 20165 43775 20223 43781
rect 20165 43741 20177 43775
rect 20211 43772 20223 43775
rect 20916 43772 20944 43948
rect 25406 43868 25412 43920
rect 25464 43908 25470 43920
rect 25777 43911 25835 43917
rect 25777 43908 25789 43911
rect 25464 43880 25789 43908
rect 25464 43868 25470 43880
rect 25777 43877 25789 43880
rect 25823 43908 25835 43911
rect 27801 43911 27859 43917
rect 25823 43880 27752 43908
rect 25823 43877 25835 43880
rect 25777 43871 25835 43877
rect 20990 43800 20996 43852
rect 21048 43840 21054 43852
rect 27341 43843 27399 43849
rect 21048 43812 22324 43840
rect 21048 43800 21054 43812
rect 20211 43744 20944 43772
rect 21085 43775 21143 43781
rect 20211 43741 20223 43744
rect 20165 43735 20223 43741
rect 21085 43741 21097 43775
rect 21131 43772 21143 43775
rect 21174 43772 21180 43784
rect 21131 43744 21180 43772
rect 21131 43741 21143 43744
rect 21085 43735 21143 43741
rect 21174 43732 21180 43744
rect 21232 43732 21238 43784
rect 21358 43772 21364 43784
rect 21319 43744 21364 43772
rect 21358 43732 21364 43744
rect 21416 43732 21422 43784
rect 21818 43772 21824 43784
rect 21468 43744 21824 43772
rect 20714 43704 20720 43716
rect 16776 43676 20720 43704
rect 20714 43664 20720 43676
rect 20772 43664 20778 43716
rect 21192 43704 21220 43732
rect 21468 43704 21496 43744
rect 21818 43732 21824 43744
rect 21876 43772 21882 43784
rect 22296 43781 22324 43812
rect 27341 43809 27353 43843
rect 27387 43809 27399 43843
rect 27724 43840 27752 43880
rect 27801 43877 27813 43911
rect 27847 43908 27859 43911
rect 27908 43908 27936 43948
rect 28994 43936 29000 43948
rect 29052 43936 29058 43988
rect 29733 43979 29791 43985
rect 29733 43945 29745 43979
rect 29779 43976 29791 43979
rect 31202 43976 31208 43988
rect 29779 43948 31208 43976
rect 29779 43945 29791 43948
rect 29733 43939 29791 43945
rect 31202 43936 31208 43948
rect 31260 43976 31266 43988
rect 34422 43976 34428 43988
rect 31260 43948 34428 43976
rect 31260 43936 31266 43948
rect 34422 43936 34428 43948
rect 34480 43936 34486 43988
rect 36354 43936 36360 43988
rect 36412 43976 36418 43988
rect 36449 43979 36507 43985
rect 36449 43976 36461 43979
rect 36412 43948 36461 43976
rect 36412 43936 36418 43948
rect 36449 43945 36461 43948
rect 36495 43945 36507 43979
rect 36449 43939 36507 43945
rect 40221 43979 40279 43985
rect 40221 43945 40233 43979
rect 40267 43976 40279 43979
rect 40402 43976 40408 43988
rect 40267 43948 40408 43976
rect 40267 43945 40279 43948
rect 40221 43939 40279 43945
rect 27847 43880 27936 43908
rect 27847 43877 27859 43880
rect 27801 43871 27859 43877
rect 28902 43868 28908 43920
rect 28960 43908 28966 43920
rect 29917 43911 29975 43917
rect 29917 43908 29929 43911
rect 28960 43880 29929 43908
rect 28960 43868 28966 43880
rect 29917 43877 29929 43880
rect 29963 43877 29975 43911
rect 29917 43871 29975 43877
rect 35802 43868 35808 43920
rect 35860 43908 35866 43920
rect 40236 43908 40264 43939
rect 40402 43936 40408 43948
rect 40460 43936 40466 43988
rect 42521 43979 42579 43985
rect 42521 43945 42533 43979
rect 42567 43976 42579 43979
rect 43162 43976 43168 43988
rect 42567 43948 43168 43976
rect 42567 43945 42579 43948
rect 42521 43939 42579 43945
rect 43162 43936 43168 43948
rect 43220 43936 43226 43988
rect 44358 43976 44364 43988
rect 44319 43948 44364 43976
rect 44358 43936 44364 43948
rect 44416 43936 44422 43988
rect 35860 43880 40264 43908
rect 35860 43868 35866 43880
rect 28194 43843 28252 43849
rect 28194 43840 28206 43843
rect 27724 43812 28206 43840
rect 27341 43803 27399 43809
rect 28194 43809 28206 43812
rect 28240 43809 28252 43843
rect 30926 43840 30932 43852
rect 30887 43812 30932 43840
rect 28194 43803 28252 43809
rect 22005 43775 22063 43781
rect 22005 43772 22017 43775
rect 21876 43744 22017 43772
rect 21876 43732 21882 43744
rect 22005 43741 22017 43744
rect 22051 43741 22063 43775
rect 22005 43735 22063 43741
rect 22281 43775 22339 43781
rect 22281 43741 22293 43775
rect 22327 43741 22339 43775
rect 22738 43772 22744 43784
rect 22699 43744 22744 43772
rect 22281 43735 22339 43741
rect 22738 43732 22744 43744
rect 22796 43732 22802 43784
rect 23017 43775 23075 43781
rect 23017 43741 23029 43775
rect 23063 43741 23075 43775
rect 23017 43735 23075 43741
rect 21910 43704 21916 43716
rect 21192 43676 21496 43704
rect 21560 43676 21916 43704
rect 21560 43648 21588 43676
rect 21910 43664 21916 43676
rect 21968 43704 21974 43716
rect 22189 43707 22247 43713
rect 22189 43704 22201 43707
rect 21968 43676 22201 43704
rect 21968 43664 21974 43676
rect 22189 43673 22201 43676
rect 22235 43704 22247 43707
rect 23032 43704 23060 43735
rect 24118 43732 24124 43784
rect 24176 43772 24182 43784
rect 24397 43775 24455 43781
rect 24397 43772 24409 43775
rect 24176 43744 24409 43772
rect 24176 43732 24182 43744
rect 24397 43741 24409 43744
rect 24443 43741 24455 43775
rect 24397 43735 24455 43741
rect 24664 43775 24722 43781
rect 24664 43741 24676 43775
rect 24710 43772 24722 43775
rect 25038 43772 25044 43784
rect 24710 43744 25044 43772
rect 24710 43741 24722 43744
rect 24664 43735 24722 43741
rect 25038 43732 25044 43744
rect 25096 43732 25102 43784
rect 26237 43775 26295 43781
rect 26237 43772 26249 43775
rect 25884 43744 26249 43772
rect 22235 43676 23060 43704
rect 22235 43673 22247 43676
rect 22189 43667 22247 43673
rect 13354 43596 13360 43648
rect 13412 43636 13418 43648
rect 13541 43639 13599 43645
rect 13541 43636 13553 43639
rect 13412 43608 13553 43636
rect 13412 43596 13418 43608
rect 13541 43605 13553 43608
rect 13587 43605 13599 43639
rect 13541 43599 13599 43605
rect 16758 43596 16764 43648
rect 16816 43636 16822 43648
rect 18141 43639 18199 43645
rect 18141 43636 18153 43639
rect 16816 43608 18153 43636
rect 16816 43596 16822 43608
rect 18141 43605 18153 43608
rect 18187 43636 18199 43639
rect 20254 43636 20260 43648
rect 18187 43608 20260 43636
rect 18187 43605 18199 43608
rect 18141 43599 18199 43605
rect 20254 43596 20260 43608
rect 20312 43596 20318 43648
rect 20901 43639 20959 43645
rect 20901 43605 20913 43639
rect 20947 43636 20959 43639
rect 21082 43636 21088 43648
rect 20947 43608 21088 43636
rect 20947 43605 20959 43608
rect 20901 43599 20959 43605
rect 21082 43596 21088 43608
rect 21140 43596 21146 43648
rect 21269 43639 21327 43645
rect 21269 43605 21281 43639
rect 21315 43636 21327 43639
rect 21542 43636 21548 43648
rect 21315 43608 21548 43636
rect 21315 43605 21327 43608
rect 21269 43599 21327 43605
rect 21542 43596 21548 43608
rect 21600 43596 21606 43648
rect 21821 43639 21879 43645
rect 21821 43605 21833 43639
rect 21867 43636 21879 43639
rect 23014 43636 23020 43648
rect 21867 43608 23020 43636
rect 21867 43605 21879 43608
rect 21821 43599 21879 43605
rect 23014 43596 23020 43608
rect 23072 43596 23078 43648
rect 24302 43596 24308 43648
rect 24360 43636 24366 43648
rect 25884 43636 25912 43744
rect 26237 43741 26249 43744
rect 26283 43741 26295 43775
rect 27154 43772 27160 43784
rect 27115 43744 27160 43772
rect 26237 43735 26295 43741
rect 27154 43732 27160 43744
rect 27212 43732 27218 43784
rect 24360 43608 25912 43636
rect 26421 43639 26479 43645
rect 24360 43596 24366 43608
rect 26421 43605 26433 43639
rect 26467 43636 26479 43639
rect 26970 43636 26976 43648
rect 26467 43608 26976 43636
rect 26467 43605 26479 43608
rect 26421 43599 26479 43605
rect 26970 43596 26976 43608
rect 27028 43596 27034 43648
rect 27356 43636 27384 43803
rect 30926 43800 30932 43812
rect 30984 43800 30990 43852
rect 34514 43800 34520 43852
rect 34572 43840 34578 43852
rect 36170 43840 36176 43852
rect 34572 43812 36176 43840
rect 34572 43800 34578 43812
rect 36170 43800 36176 43812
rect 36228 43840 36234 43852
rect 36541 43843 36599 43849
rect 36541 43840 36553 43843
rect 36228 43812 36553 43840
rect 36228 43800 36234 43812
rect 36541 43809 36553 43812
rect 36587 43809 36599 43843
rect 36541 43803 36599 43809
rect 38654 43800 38660 43852
rect 38712 43840 38718 43852
rect 38838 43840 38844 43852
rect 38712 43812 38844 43840
rect 38712 43800 38718 43812
rect 38838 43800 38844 43812
rect 38896 43800 38902 43852
rect 43993 43843 44051 43849
rect 43993 43809 44005 43843
rect 44039 43840 44051 43843
rect 44910 43840 44916 43852
rect 44039 43812 44916 43840
rect 44039 43809 44051 43812
rect 43993 43803 44051 43809
rect 44910 43800 44916 43812
rect 44968 43800 44974 43852
rect 45646 43840 45652 43852
rect 45607 43812 45652 43840
rect 45646 43800 45652 43812
rect 45704 43800 45710 43852
rect 66257 43843 66315 43849
rect 66257 43809 66269 43843
rect 66303 43840 66315 43843
rect 67910 43840 67916 43852
rect 66303 43812 67916 43840
rect 66303 43809 66315 43812
rect 66257 43803 66315 43809
rect 67910 43800 67916 43812
rect 67968 43800 67974 43852
rect 28074 43732 28080 43784
rect 28132 43772 28138 43784
rect 28350 43772 28356 43784
rect 28132 43744 28177 43772
rect 28311 43744 28356 43772
rect 28132 43732 28138 43744
rect 28350 43732 28356 43744
rect 28408 43732 28414 43784
rect 28997 43775 29055 43781
rect 28997 43741 29009 43775
rect 29043 43772 29055 43775
rect 31196 43775 31254 43781
rect 29043 43744 31156 43772
rect 29043 43741 29055 43744
rect 28997 43735 29055 43741
rect 29546 43704 29552 43716
rect 29507 43676 29552 43704
rect 29546 43664 29552 43676
rect 29604 43664 29610 43716
rect 29765 43707 29823 43713
rect 29765 43673 29777 43707
rect 29811 43704 29823 43707
rect 29914 43704 29920 43716
rect 29811 43676 29920 43704
rect 29811 43673 29823 43676
rect 29765 43667 29823 43673
rect 29914 43664 29920 43676
rect 29972 43664 29978 43716
rect 31128 43704 31156 43744
rect 31196 43741 31208 43775
rect 31242 43772 31254 43775
rect 32122 43772 32128 43784
rect 31242 43744 32128 43772
rect 31242 43741 31254 43744
rect 31196 43735 31254 43741
rect 32122 43732 32128 43744
rect 32180 43732 32186 43784
rect 32766 43772 32772 43784
rect 32727 43744 32772 43772
rect 32766 43732 32772 43744
rect 32824 43732 32830 43784
rect 33036 43775 33094 43781
rect 33036 43741 33048 43775
rect 33082 43772 33094 43775
rect 33778 43772 33784 43784
rect 33082 43744 33784 43772
rect 33082 43741 33094 43744
rect 33036 43735 33094 43741
rect 33778 43732 33784 43744
rect 33836 43732 33842 43784
rect 36262 43772 36268 43784
rect 36223 43744 36268 43772
rect 36262 43732 36268 43744
rect 36320 43732 36326 43784
rect 37918 43772 37924 43784
rect 37879 43744 37924 43772
rect 37918 43732 37924 43744
rect 37976 43732 37982 43784
rect 38102 43772 38108 43784
rect 38063 43744 38108 43772
rect 38102 43732 38108 43744
rect 38160 43732 38166 43784
rect 38197 43775 38255 43781
rect 38197 43741 38209 43775
rect 38243 43772 38255 43775
rect 38930 43772 38936 43784
rect 38243 43744 38936 43772
rect 38243 43741 38255 43744
rect 38197 43735 38255 43741
rect 38930 43732 38936 43744
rect 38988 43732 38994 43784
rect 40037 43775 40095 43781
rect 40037 43741 40049 43775
rect 40083 43772 40095 43775
rect 40494 43772 40500 43784
rect 40083 43744 40500 43772
rect 40083 43741 40095 43744
rect 40037 43735 40095 43741
rect 40494 43732 40500 43744
rect 40552 43772 40558 43784
rect 40865 43775 40923 43781
rect 40865 43772 40877 43775
rect 40552 43744 40877 43772
rect 40552 43732 40558 43744
rect 40865 43741 40877 43744
rect 40911 43741 40923 43775
rect 42426 43772 42432 43784
rect 42387 43744 42432 43772
rect 40865 43735 40923 43741
rect 42426 43732 42432 43744
rect 42484 43732 42490 43784
rect 44174 43772 44180 43784
rect 44135 43744 44180 43772
rect 44174 43732 44180 43744
rect 44232 43732 44238 43784
rect 46198 43732 46204 43784
rect 46256 43772 46262 43784
rect 48041 43775 48099 43781
rect 46256 43744 47716 43772
rect 46256 43732 46262 43744
rect 35986 43704 35992 43716
rect 31128 43676 35992 43704
rect 35986 43664 35992 43676
rect 36044 43664 36050 43716
rect 36081 43707 36139 43713
rect 36081 43673 36093 43707
rect 36127 43704 36139 43707
rect 38120 43704 38148 43732
rect 38654 43704 38660 43716
rect 36127 43676 38148 43704
rect 38615 43676 38660 43704
rect 36127 43673 36139 43676
rect 36081 43667 36139 43673
rect 38654 43664 38660 43676
rect 38712 43664 38718 43716
rect 38838 43704 38844 43716
rect 38799 43676 38844 43704
rect 38838 43664 38844 43676
rect 38896 43664 38902 43716
rect 41049 43707 41107 43713
rect 41049 43673 41061 43707
rect 41095 43704 41107 43707
rect 42518 43704 42524 43716
rect 41095 43676 42524 43704
rect 41095 43673 41107 43676
rect 41049 43667 41107 43673
rect 42518 43664 42524 43676
rect 42576 43664 42582 43716
rect 45916 43707 45974 43713
rect 45916 43673 45928 43707
rect 45962 43704 45974 43707
rect 46382 43704 46388 43716
rect 45962 43676 46388 43704
rect 45962 43673 45974 43676
rect 45916 43667 45974 43673
rect 46382 43664 46388 43676
rect 46440 43664 46446 43716
rect 47688 43648 47716 43744
rect 48041 43741 48053 43775
rect 48087 43772 48099 43775
rect 48590 43772 48596 43784
rect 48087 43744 48596 43772
rect 48087 43741 48099 43744
rect 48041 43735 48099 43741
rect 48590 43732 48596 43744
rect 48648 43732 48654 43784
rect 48314 43713 48320 43716
rect 48308 43667 48320 43713
rect 48372 43704 48378 43716
rect 66438 43704 66444 43716
rect 48372 43676 48408 43704
rect 66399 43676 66444 43704
rect 48314 43664 48320 43667
rect 48372 43664 48378 43676
rect 66438 43664 66444 43676
rect 66496 43664 66502 43716
rect 68094 43704 68100 43716
rect 68055 43676 68100 43704
rect 68094 43664 68100 43676
rect 68152 43664 68158 43716
rect 28810 43636 28816 43648
rect 27356 43608 28816 43636
rect 28810 43596 28816 43608
rect 28868 43596 28874 43648
rect 30742 43596 30748 43648
rect 30800 43636 30806 43648
rect 32309 43639 32367 43645
rect 32309 43636 32321 43639
rect 30800 43608 32321 43636
rect 30800 43596 30806 43608
rect 32309 43605 32321 43608
rect 32355 43605 32367 43639
rect 32309 43599 32367 43605
rect 33594 43596 33600 43648
rect 33652 43636 33658 43648
rect 34149 43639 34207 43645
rect 34149 43636 34161 43639
rect 33652 43608 34161 43636
rect 33652 43596 33658 43608
rect 34149 43605 34161 43608
rect 34195 43605 34207 43639
rect 34149 43599 34207 43605
rect 38470 43596 38476 43648
rect 38528 43636 38534 43648
rect 39025 43639 39083 43645
rect 39025 43636 39037 43639
rect 38528 43608 39037 43636
rect 38528 43596 38534 43608
rect 39025 43605 39037 43608
rect 39071 43605 39083 43639
rect 39025 43599 39083 43605
rect 45646 43596 45652 43648
rect 45704 43636 45710 43648
rect 47029 43639 47087 43645
rect 47029 43636 47041 43639
rect 45704 43608 47041 43636
rect 45704 43596 45710 43608
rect 47029 43605 47041 43608
rect 47075 43605 47087 43639
rect 47029 43599 47087 43605
rect 47670 43596 47676 43648
rect 47728 43636 47734 43648
rect 49421 43639 49479 43645
rect 49421 43636 49433 43639
rect 47728 43608 49433 43636
rect 47728 43596 47734 43608
rect 49421 43605 49433 43608
rect 49467 43605 49479 43639
rect 49421 43599 49479 43605
rect 1104 43546 68816 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 68816 43546
rect 1104 43472 68816 43494
rect 14642 43392 14648 43444
rect 14700 43432 14706 43444
rect 14737 43435 14795 43441
rect 14737 43432 14749 43435
rect 14700 43404 14749 43432
rect 14700 43392 14706 43404
rect 14737 43401 14749 43404
rect 14783 43401 14795 43435
rect 14737 43395 14795 43401
rect 15378 43392 15384 43444
rect 15436 43432 15442 43444
rect 15657 43435 15715 43441
rect 15657 43432 15669 43435
rect 15436 43404 15669 43432
rect 15436 43392 15442 43404
rect 15657 43401 15669 43404
rect 15703 43401 15715 43435
rect 15657 43395 15715 43401
rect 15746 43392 15752 43444
rect 15804 43432 15810 43444
rect 17034 43432 17040 43444
rect 15804 43404 16896 43432
rect 16995 43404 17040 43432
rect 15804 43392 15810 43404
rect 16574 43364 16580 43376
rect 15396 43336 16580 43364
rect 12618 43256 12624 43308
rect 12676 43296 12682 43308
rect 12986 43305 12992 43308
rect 12713 43299 12771 43305
rect 12713 43296 12725 43299
rect 12676 43268 12725 43296
rect 12676 43256 12682 43268
rect 12713 43265 12725 43268
rect 12759 43265 12771 43299
rect 12713 43259 12771 43265
rect 12980 43259 12992 43305
rect 13044 43296 13050 43308
rect 14550 43296 14556 43308
rect 13044 43268 13080 43296
rect 14511 43268 14556 43296
rect 12986 43256 12992 43259
rect 13044 43256 13050 43268
rect 14550 43256 14556 43268
rect 14608 43256 14614 43308
rect 15396 43305 15424 43336
rect 16574 43324 16580 43336
rect 16632 43324 16638 43376
rect 15381 43299 15439 43305
rect 15381 43265 15393 43299
rect 15427 43265 15439 43299
rect 15381 43259 15439 43265
rect 15473 43299 15531 43305
rect 15473 43265 15485 43299
rect 15519 43296 15531 43299
rect 15562 43296 15568 43308
rect 15519 43268 15568 43296
rect 15519 43265 15531 43268
rect 15473 43259 15531 43265
rect 15562 43256 15568 43268
rect 15620 43256 15626 43308
rect 16758 43296 16764 43308
rect 16719 43268 16764 43296
rect 16758 43256 16764 43268
rect 16816 43256 16822 43308
rect 16868 43305 16896 43404
rect 17034 43392 17040 43404
rect 17092 43392 17098 43444
rect 19150 43392 19156 43444
rect 19208 43432 19214 43444
rect 20438 43432 20444 43444
rect 19208 43404 20444 43432
rect 19208 43392 19214 43404
rect 20438 43392 20444 43404
rect 20496 43392 20502 43444
rect 20530 43392 20536 43444
rect 20588 43432 20594 43444
rect 24118 43432 24124 43444
rect 20588 43404 23980 43432
rect 24079 43404 24124 43432
rect 20588 43392 20594 43404
rect 23952 43364 23980 43404
rect 24118 43392 24124 43404
rect 24176 43392 24182 43444
rect 25222 43392 25228 43444
rect 25280 43432 25286 43444
rect 25685 43435 25743 43441
rect 25685 43432 25697 43435
rect 25280 43404 25697 43432
rect 25280 43392 25286 43404
rect 25685 43401 25697 43404
rect 25731 43401 25743 43435
rect 25685 43395 25743 43401
rect 27154 43392 27160 43444
rect 27212 43432 27218 43444
rect 28353 43435 28411 43441
rect 28353 43432 28365 43435
rect 27212 43404 28365 43432
rect 27212 43392 27218 43404
rect 28353 43401 28365 43404
rect 28399 43432 28411 43435
rect 29546 43432 29552 43444
rect 28399 43404 29552 43432
rect 28399 43401 28411 43404
rect 28353 43395 28411 43401
rect 29546 43392 29552 43404
rect 29604 43392 29610 43444
rect 29638 43392 29644 43444
rect 29696 43432 29702 43444
rect 30466 43432 30472 43444
rect 29696 43404 30472 43432
rect 29696 43392 29702 43404
rect 30466 43392 30472 43404
rect 30524 43392 30530 43444
rect 32766 43392 32772 43444
rect 32824 43432 32830 43444
rect 33229 43435 33287 43441
rect 33229 43432 33241 43435
rect 32824 43404 33241 43432
rect 32824 43392 32830 43404
rect 33229 43401 33241 43404
rect 33275 43401 33287 43435
rect 34146 43432 34152 43444
rect 34107 43404 34152 43432
rect 33229 43395 33287 43401
rect 34146 43392 34152 43404
rect 34204 43392 34210 43444
rect 38838 43392 38844 43444
rect 38896 43432 38902 43444
rect 39850 43432 39856 43444
rect 38896 43404 39856 43432
rect 38896 43392 38902 43404
rect 39850 43392 39856 43404
rect 39908 43432 39914 43444
rect 40221 43435 40279 43441
rect 40221 43432 40233 43435
rect 39908 43404 40233 43432
rect 39908 43392 39914 43404
rect 40221 43401 40233 43404
rect 40267 43401 40279 43435
rect 46382 43432 46388 43444
rect 46343 43404 46388 43432
rect 40221 43395 40279 43401
rect 46382 43392 46388 43404
rect 46440 43392 46446 43444
rect 48498 43392 48504 43444
rect 48556 43432 48562 43444
rect 48593 43435 48651 43441
rect 48593 43432 48605 43435
rect 48556 43404 48605 43432
rect 48556 43392 48562 43404
rect 48593 43401 48605 43404
rect 48639 43401 48651 43435
rect 48593 43395 48651 43401
rect 66438 43392 66444 43444
rect 66496 43432 66502 43444
rect 67545 43435 67603 43441
rect 67545 43432 67557 43435
rect 66496 43404 67557 43432
rect 66496 43392 66502 43404
rect 67545 43401 67557 43404
rect 67591 43401 67603 43435
rect 67545 43395 67603 43401
rect 25774 43364 25780 43376
rect 23952 43336 25780 43364
rect 25774 43324 25780 43336
rect 25832 43324 25838 43376
rect 27246 43373 27252 43376
rect 27240 43364 27252 43373
rect 27207 43336 27252 43364
rect 27240 43327 27252 43336
rect 27246 43324 27252 43327
rect 27304 43324 27310 43376
rect 33594 43324 33600 43376
rect 33652 43364 33658 43376
rect 33781 43367 33839 43373
rect 33781 43364 33793 43367
rect 33652 43336 33793 43364
rect 33652 43324 33658 43336
rect 33781 43333 33793 43336
rect 33827 43333 33839 43367
rect 33781 43327 33839 43333
rect 33962 43324 33968 43376
rect 34020 43373 34026 43376
rect 34020 43367 34039 43373
rect 34027 43333 34039 43367
rect 34020 43327 34039 43333
rect 34020 43324 34026 43327
rect 34514 43324 34520 43376
rect 34572 43364 34578 43376
rect 34701 43367 34759 43373
rect 34701 43364 34713 43367
rect 34572 43336 34713 43364
rect 34572 43324 34578 43336
rect 34701 43333 34713 43336
rect 34747 43333 34759 43367
rect 34701 43327 34759 43333
rect 38381 43367 38439 43373
rect 38381 43333 38393 43367
rect 38427 43364 38439 43367
rect 38654 43364 38660 43376
rect 38427 43336 38660 43364
rect 38427 43333 38439 43336
rect 38381 43327 38439 43333
rect 16853 43299 16911 43305
rect 16853 43265 16865 43299
rect 16899 43265 16911 43299
rect 16853 43259 16911 43265
rect 20254 43256 20260 43308
rect 20312 43305 20318 43308
rect 20312 43299 20340 43305
rect 20328 43265 20340 43299
rect 22554 43296 22560 43308
rect 22515 43268 22560 43296
rect 20312 43259 20340 43265
rect 20312 43256 20318 43259
rect 22554 43256 22560 43268
rect 22612 43256 22618 43308
rect 24026 43296 24032 43308
rect 23987 43268 24032 43296
rect 24026 43256 24032 43268
rect 24084 43256 24090 43308
rect 25406 43296 25412 43308
rect 25367 43268 25412 43296
rect 25406 43256 25412 43268
rect 25464 43256 25470 43308
rect 25501 43299 25559 43305
rect 25501 43265 25513 43299
rect 25547 43265 25559 43299
rect 26970 43296 26976 43308
rect 26931 43268 26976 43296
rect 25501 43259 25559 43265
rect 19245 43231 19303 43237
rect 19245 43197 19257 43231
rect 19291 43228 19303 43231
rect 19334 43228 19340 43240
rect 19291 43200 19340 43228
rect 19291 43197 19303 43200
rect 19245 43191 19303 43197
rect 19334 43188 19340 43200
rect 19392 43188 19398 43240
rect 19429 43231 19487 43237
rect 19429 43197 19441 43231
rect 19475 43228 19487 43231
rect 20162 43228 20168 43240
rect 19475 43200 20024 43228
rect 20123 43200 20168 43228
rect 19475 43197 19487 43200
rect 19429 43191 19487 43197
rect 14090 43160 14096 43172
rect 14003 43132 14096 43160
rect 14090 43120 14096 43132
rect 14148 43160 14154 43172
rect 18966 43160 18972 43172
rect 14148 43132 18972 43160
rect 14148 43120 14154 43132
rect 18966 43120 18972 43132
rect 19024 43120 19030 43172
rect 19058 43120 19064 43172
rect 19116 43160 19122 43172
rect 19889 43163 19947 43169
rect 19889 43160 19901 43163
rect 19116 43132 19901 43160
rect 19116 43120 19122 43132
rect 19889 43129 19901 43132
rect 19935 43129 19947 43163
rect 19889 43123 19947 43129
rect 19996 43092 20024 43200
rect 20162 43188 20168 43200
rect 20220 43188 20226 43240
rect 20438 43228 20444 43240
rect 20399 43200 20444 43228
rect 20438 43188 20444 43200
rect 20496 43188 20502 43240
rect 21174 43188 21180 43240
rect 21232 43228 21238 43240
rect 22833 43231 22891 43237
rect 22833 43228 22845 43231
rect 21232 43200 22845 43228
rect 21232 43188 21238 43200
rect 22833 43197 22845 43200
rect 22879 43197 22891 43231
rect 22833 43191 22891 43197
rect 25222 43188 25228 43240
rect 25280 43228 25286 43240
rect 25516 43228 25544 43259
rect 26970 43256 26976 43268
rect 27028 43256 27034 43308
rect 28994 43256 29000 43308
rect 29052 43296 29058 43308
rect 29365 43299 29423 43305
rect 29052 43268 29316 43296
rect 29052 43256 29058 43268
rect 25280 43200 25544 43228
rect 29181 43231 29239 43237
rect 25280 43188 25286 43200
rect 29181 43197 29193 43231
rect 29227 43197 29239 43231
rect 29181 43191 29239 43197
rect 21266 43160 21272 43172
rect 21008 43132 21272 43160
rect 21008 43092 21036 43132
rect 21266 43120 21272 43132
rect 21324 43120 21330 43172
rect 19996 43064 21036 43092
rect 21085 43095 21143 43101
rect 21085 43061 21097 43095
rect 21131 43092 21143 43095
rect 21634 43092 21640 43104
rect 21131 43064 21640 43092
rect 21131 43061 21143 43064
rect 21085 43055 21143 43061
rect 21634 43052 21640 43064
rect 21692 43052 21698 43104
rect 29196 43092 29224 43191
rect 29288 43160 29316 43268
rect 29365 43265 29377 43299
rect 29411 43296 29423 43299
rect 29546 43296 29552 43308
rect 29411 43268 29552 43296
rect 29411 43265 29423 43268
rect 29365 43259 29423 43265
rect 29546 43256 29552 43268
rect 29604 43256 29610 43308
rect 33229 43299 33287 43305
rect 33229 43265 33241 43299
rect 33275 43296 33287 43299
rect 33870 43296 33876 43308
rect 33275 43268 33876 43296
rect 33275 43265 33287 43268
rect 33229 43259 33287 43265
rect 33870 43256 33876 43268
rect 33928 43256 33934 43308
rect 37826 43256 37832 43308
rect 37884 43296 37890 43308
rect 38013 43299 38071 43305
rect 38013 43296 38025 43299
rect 37884 43268 38025 43296
rect 37884 43256 37890 43268
rect 38013 43265 38025 43268
rect 38059 43265 38071 43299
rect 38013 43259 38071 43265
rect 29454 43188 29460 43240
rect 29512 43228 29518 43240
rect 30101 43231 30159 43237
rect 30101 43228 30113 43231
rect 29512 43200 30113 43228
rect 29512 43188 29518 43200
rect 30101 43197 30113 43200
rect 30147 43197 30159 43231
rect 30101 43191 30159 43197
rect 30190 43188 30196 43240
rect 30248 43237 30254 43240
rect 30248 43231 30276 43237
rect 30264 43197 30276 43231
rect 30248 43191 30276 43197
rect 30377 43231 30435 43237
rect 30377 43197 30389 43231
rect 30423 43228 30435 43231
rect 30558 43228 30564 43240
rect 30423 43200 30564 43228
rect 30423 43197 30435 43200
rect 30377 43191 30435 43197
rect 30248 43188 30254 43191
rect 30558 43188 30564 43200
rect 30616 43188 30622 43240
rect 31018 43188 31024 43240
rect 31076 43228 31082 43240
rect 38396 43228 38424 43327
rect 38654 43324 38660 43336
rect 38712 43324 38718 43376
rect 40494 43324 40500 43376
rect 40552 43364 40558 43376
rect 40773 43367 40831 43373
rect 40773 43364 40785 43367
rect 40552 43336 40785 43364
rect 40552 43324 40558 43336
rect 40773 43333 40785 43336
rect 40819 43333 40831 43367
rect 40773 43327 40831 43333
rect 44008 43336 48452 43364
rect 39108 43299 39166 43305
rect 39108 43265 39120 43299
rect 39154 43296 39166 43299
rect 39390 43296 39396 43308
rect 39154 43268 39396 43296
rect 39154 43265 39166 43268
rect 39108 43259 39166 43265
rect 39390 43256 39396 43268
rect 39448 43256 39454 43308
rect 41785 43299 41843 43305
rect 41785 43265 41797 43299
rect 41831 43296 41843 43299
rect 42518 43296 42524 43308
rect 41831 43268 42524 43296
rect 41831 43265 41843 43268
rect 41785 43259 41843 43265
rect 42518 43256 42524 43268
rect 42576 43296 42582 43308
rect 44008 43305 44036 43336
rect 43993 43299 44051 43305
rect 43993 43296 44005 43299
rect 42576 43268 44005 43296
rect 42576 43256 42582 43268
rect 43993 43265 44005 43268
rect 44039 43265 44051 43299
rect 45646 43296 45652 43308
rect 45607 43268 45652 43296
rect 43993 43259 44051 43265
rect 45646 43256 45652 43268
rect 45704 43256 45710 43308
rect 45741 43299 45799 43305
rect 45741 43265 45753 43299
rect 45787 43265 45799 43299
rect 45741 43259 45799 43265
rect 45925 43299 45983 43305
rect 45925 43265 45937 43299
rect 45971 43296 45983 43299
rect 46569 43299 46627 43305
rect 46569 43296 46581 43299
rect 45971 43268 46581 43296
rect 45971 43265 45983 43268
rect 45925 43259 45983 43265
rect 46569 43265 46581 43268
rect 46615 43265 46627 43299
rect 47670 43296 47676 43308
rect 47631 43268 47676 43296
rect 46569 43259 46627 43265
rect 38838 43228 38844 43240
rect 31076 43200 38424 43228
rect 38799 43200 38844 43228
rect 31076 43188 31082 43200
rect 38838 43188 38844 43200
rect 38896 43188 38902 43240
rect 44174 43188 44180 43240
rect 44232 43228 44238 43240
rect 45756 43228 45784 43259
rect 47670 43256 47676 43268
rect 47728 43256 47734 43308
rect 47762 43256 47768 43308
rect 47820 43296 47826 43308
rect 48424 43305 48452 43336
rect 48409 43299 48467 43305
rect 47820 43268 47913 43296
rect 47820 43256 47826 43268
rect 48409 43265 48421 43299
rect 48455 43296 48467 43299
rect 48682 43296 48688 43308
rect 48455 43268 48688 43296
rect 48455 43265 48467 43268
rect 48409 43259 48467 43265
rect 48682 43256 48688 43268
rect 48740 43256 48746 43308
rect 66990 43256 66996 43308
rect 67048 43296 67054 43308
rect 67453 43299 67511 43305
rect 67453 43296 67465 43299
rect 67048 43268 67465 43296
rect 67048 43256 67054 43268
rect 67453 43265 67465 43268
rect 67499 43265 67511 43299
rect 67453 43259 67511 43265
rect 47780 43228 47808 43256
rect 44232 43200 47808 43228
rect 44232 43188 44238 43200
rect 29825 43163 29883 43169
rect 29825 43160 29837 43163
rect 29288 43132 29837 43160
rect 29825 43129 29837 43132
rect 29871 43129 29883 43163
rect 29825 43123 29883 43129
rect 31754 43120 31760 43172
rect 31812 43160 31818 43172
rect 35894 43160 35900 43172
rect 31812 43132 35900 43160
rect 31812 43120 31818 43132
rect 35894 43120 35900 43132
rect 35952 43120 35958 43172
rect 40954 43160 40960 43172
rect 40915 43132 40960 43160
rect 40954 43120 40960 43132
rect 41012 43120 41018 43172
rect 30742 43092 30748 43104
rect 29196 43064 30748 43092
rect 30742 43052 30748 43064
rect 30800 43052 30806 43104
rect 31021 43095 31079 43101
rect 31021 43061 31033 43095
rect 31067 43092 31079 43095
rect 32950 43092 32956 43104
rect 31067 43064 32956 43092
rect 31067 43061 31079 43064
rect 31021 43055 31079 43061
rect 32950 43052 32956 43064
rect 33008 43052 33014 43104
rect 33965 43095 34023 43101
rect 33965 43061 33977 43095
rect 34011 43092 34023 43095
rect 34422 43092 34428 43104
rect 34011 43064 34428 43092
rect 34011 43061 34023 43064
rect 33965 43055 34023 43061
rect 34422 43052 34428 43064
rect 34480 43052 34486 43104
rect 34514 43052 34520 43104
rect 34572 43092 34578 43104
rect 34793 43095 34851 43101
rect 34793 43092 34805 43095
rect 34572 43064 34805 43092
rect 34572 43052 34578 43064
rect 34793 43061 34805 43064
rect 34839 43061 34851 43095
rect 41782 43092 41788 43104
rect 41743 43064 41788 43092
rect 34793 43055 34851 43061
rect 41782 43052 41788 43064
rect 41840 43052 41846 43104
rect 43806 43092 43812 43104
rect 43767 43064 43812 43092
rect 43806 43052 43812 43064
rect 43864 43052 43870 43104
rect 47949 43095 48007 43101
rect 47949 43061 47961 43095
rect 47995 43092 48007 43095
rect 48130 43092 48136 43104
rect 47995 43064 48136 43092
rect 47995 43061 48007 43064
rect 47949 43055 48007 43061
rect 48130 43052 48136 43064
rect 48188 43052 48194 43104
rect 1104 43002 68816 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 65654 43002
rect 65706 42950 65718 43002
rect 65770 42950 65782 43002
rect 65834 42950 65846 43002
rect 65898 42950 65910 43002
rect 65962 42950 68816 43002
rect 1104 42928 68816 42950
rect 12986 42848 12992 42900
rect 13044 42888 13050 42900
rect 13173 42891 13231 42897
rect 13173 42888 13185 42891
rect 13044 42860 13185 42888
rect 13044 42848 13050 42860
rect 13173 42857 13185 42860
rect 13219 42857 13231 42891
rect 13173 42851 13231 42857
rect 22738 42848 22744 42900
rect 22796 42888 22802 42900
rect 31018 42888 31024 42900
rect 22796 42860 31024 42888
rect 22796 42848 22802 42860
rect 31018 42848 31024 42860
rect 31076 42848 31082 42900
rect 32585 42891 32643 42897
rect 32585 42857 32597 42891
rect 32631 42888 32643 42891
rect 33965 42891 34023 42897
rect 33965 42888 33977 42891
rect 32631 42860 33977 42888
rect 32631 42857 32643 42860
rect 32585 42851 32643 42857
rect 33965 42857 33977 42860
rect 34011 42888 34023 42891
rect 34422 42888 34428 42900
rect 34011 42860 34428 42888
rect 34011 42857 34023 42860
rect 33965 42851 34023 42857
rect 34422 42848 34428 42860
rect 34480 42848 34486 42900
rect 38838 42848 38844 42900
rect 38896 42888 38902 42900
rect 38933 42891 38991 42897
rect 38933 42888 38945 42891
rect 38896 42860 38945 42888
rect 38896 42848 38902 42860
rect 38933 42857 38945 42860
rect 38979 42857 38991 42891
rect 38933 42851 38991 42857
rect 39942 42848 39948 42900
rect 40000 42888 40006 42900
rect 40000 42860 44220 42888
rect 40000 42848 40006 42860
rect 32766 42820 32772 42832
rect 32727 42792 32772 42820
rect 32766 42780 32772 42792
rect 32824 42780 32830 42832
rect 17589 42755 17647 42761
rect 17589 42721 17601 42755
rect 17635 42752 17647 42755
rect 17954 42752 17960 42764
rect 17635 42724 17960 42752
rect 17635 42721 17647 42724
rect 17589 42715 17647 42721
rect 17954 42712 17960 42724
rect 18012 42712 18018 42764
rect 21174 42712 21180 42764
rect 21232 42752 21238 42764
rect 21232 42724 21404 42752
rect 21232 42712 21238 42724
rect 13354 42684 13360 42696
rect 13315 42656 13360 42684
rect 13354 42644 13360 42656
rect 13412 42644 13418 42696
rect 14550 42644 14556 42696
rect 14608 42684 14614 42696
rect 14737 42687 14795 42693
rect 14737 42684 14749 42687
rect 14608 42656 14749 42684
rect 14608 42644 14614 42656
rect 14737 42653 14749 42656
rect 14783 42653 14795 42687
rect 14737 42647 14795 42653
rect 15657 42687 15715 42693
rect 15657 42653 15669 42687
rect 15703 42684 15715 42687
rect 15746 42684 15752 42696
rect 15703 42656 15752 42684
rect 15703 42653 15715 42656
rect 15657 42647 15715 42653
rect 15746 42644 15752 42656
rect 15804 42644 15810 42696
rect 16942 42684 16948 42696
rect 16903 42656 16948 42684
rect 16942 42644 16948 42656
rect 17000 42644 17006 42696
rect 17494 42644 17500 42696
rect 17552 42684 17558 42696
rect 21376 42693 21404 42724
rect 25682 42712 25688 42764
rect 25740 42752 25746 42764
rect 26050 42752 26056 42764
rect 25740 42724 26056 42752
rect 25740 42712 25746 42724
rect 26050 42712 26056 42724
rect 26108 42712 26114 42764
rect 28350 42712 28356 42764
rect 28408 42752 28414 42764
rect 31754 42752 31760 42764
rect 28408 42724 31760 42752
rect 28408 42712 28414 42724
rect 31754 42712 31760 42724
rect 31812 42712 31818 42764
rect 36262 42712 36268 42764
rect 36320 42752 36326 42764
rect 36817 42755 36875 42761
rect 36817 42752 36829 42755
rect 36320 42724 36829 42752
rect 36320 42712 36326 42724
rect 36817 42721 36829 42724
rect 36863 42752 36875 42755
rect 39850 42752 39856 42764
rect 36863 42724 38332 42752
rect 39811 42724 39856 42752
rect 36863 42721 36875 42724
rect 36817 42715 36875 42721
rect 17773 42687 17831 42693
rect 17773 42684 17785 42687
rect 17552 42656 17785 42684
rect 17552 42644 17558 42656
rect 17773 42653 17785 42656
rect 17819 42653 17831 42687
rect 17773 42647 17831 42653
rect 21361 42687 21419 42693
rect 21361 42653 21373 42687
rect 21407 42653 21419 42687
rect 21634 42684 21640 42696
rect 21595 42656 21640 42684
rect 21361 42647 21419 42653
rect 21634 42644 21640 42656
rect 21692 42644 21698 42696
rect 23661 42687 23719 42693
rect 23661 42653 23673 42687
rect 23707 42653 23719 42687
rect 23661 42647 23719 42653
rect 23753 42687 23811 42693
rect 23753 42653 23765 42687
rect 23799 42684 23811 42687
rect 24397 42687 24455 42693
rect 24397 42684 24409 42687
rect 23799 42656 24409 42684
rect 23799 42653 23811 42656
rect 23753 42647 23811 42653
rect 24397 42653 24409 42656
rect 24443 42653 24455 42687
rect 24397 42647 24455 42653
rect 1854 42616 1860 42628
rect 1815 42588 1860 42616
rect 1854 42576 1860 42588
rect 1912 42576 1918 42628
rect 16960 42616 16988 42644
rect 18782 42616 18788 42628
rect 16960 42588 18788 42616
rect 18782 42576 18788 42588
rect 18840 42616 18846 42628
rect 20990 42616 20996 42628
rect 18840 42588 20996 42616
rect 18840 42576 18846 42588
rect 20990 42576 20996 42588
rect 21048 42576 21054 42628
rect 21177 42619 21235 42625
rect 21177 42585 21189 42619
rect 21223 42616 21235 42619
rect 22278 42616 22284 42628
rect 21223 42588 22284 42616
rect 21223 42585 21235 42588
rect 21177 42579 21235 42585
rect 22278 42576 22284 42588
rect 22336 42576 22342 42628
rect 23676 42616 23704 42647
rect 25038 42644 25044 42696
rect 25096 42684 25102 42696
rect 26970 42684 26976 42696
rect 25096 42656 26976 42684
rect 25096 42644 25102 42656
rect 26970 42644 26976 42656
rect 27028 42644 27034 42696
rect 29546 42684 29552 42696
rect 29507 42656 29552 42684
rect 29546 42644 29552 42656
rect 29604 42644 29610 42696
rect 29825 42687 29883 42693
rect 29825 42653 29837 42687
rect 29871 42653 29883 42687
rect 29825 42647 29883 42653
rect 24026 42616 24032 42628
rect 23676 42588 24032 42616
rect 24026 42576 24032 42588
rect 24084 42576 24090 42628
rect 24486 42576 24492 42628
rect 24544 42616 24550 42628
rect 24642 42619 24700 42625
rect 24642 42616 24654 42619
rect 24544 42588 24654 42616
rect 24544 42576 24550 42588
rect 24642 42585 24654 42588
rect 24688 42585 24700 42619
rect 29730 42616 29736 42628
rect 24642 42579 24700 42585
rect 24780 42588 29736 42616
rect 1946 42548 1952 42560
rect 1907 42520 1952 42548
rect 1946 42508 1952 42520
rect 2004 42508 2010 42560
rect 14734 42508 14740 42560
rect 14792 42548 14798 42560
rect 14921 42551 14979 42557
rect 14921 42548 14933 42551
rect 14792 42520 14933 42548
rect 14792 42508 14798 42520
rect 14921 42517 14933 42520
rect 14967 42517 14979 42551
rect 15470 42548 15476 42560
rect 15431 42520 15476 42548
rect 14921 42511 14979 42517
rect 15470 42508 15476 42520
rect 15528 42508 15534 42560
rect 16942 42508 16948 42560
rect 17000 42548 17006 42560
rect 17037 42551 17095 42557
rect 17037 42548 17049 42551
rect 17000 42520 17049 42548
rect 17000 42508 17006 42520
rect 17037 42517 17049 42520
rect 17083 42517 17095 42551
rect 17954 42548 17960 42560
rect 17915 42520 17960 42548
rect 17037 42511 17095 42517
rect 17954 42508 17960 42520
rect 18012 42508 18018 42560
rect 21542 42548 21548 42560
rect 21503 42520 21548 42548
rect 21542 42508 21548 42520
rect 21600 42508 21606 42560
rect 23658 42508 23664 42560
rect 23716 42548 23722 42560
rect 24780 42548 24808 42588
rect 29730 42576 29736 42588
rect 29788 42576 29794 42628
rect 29840 42616 29868 42647
rect 30742 42644 30748 42696
rect 30800 42684 30806 42696
rect 30837 42687 30895 42693
rect 30837 42684 30849 42687
rect 30800 42656 30849 42684
rect 30800 42644 30806 42656
rect 30837 42653 30849 42656
rect 30883 42653 30895 42687
rect 30837 42647 30895 42653
rect 31941 42687 31999 42693
rect 31941 42653 31953 42687
rect 31987 42684 31999 42687
rect 32766 42684 32772 42696
rect 31987 42656 32772 42684
rect 31987 42653 31999 42656
rect 31941 42647 31999 42653
rect 32766 42644 32772 42656
rect 32824 42644 32830 42696
rect 34146 42644 34152 42696
rect 34204 42684 34210 42696
rect 34701 42687 34759 42693
rect 34701 42684 34713 42687
rect 34204 42656 34713 42684
rect 34204 42644 34210 42656
rect 34701 42653 34713 42656
rect 34747 42653 34759 42687
rect 34701 42647 34759 42653
rect 37093 42687 37151 42693
rect 37093 42653 37105 42687
rect 37139 42684 37151 42687
rect 37366 42684 37372 42696
rect 37139 42656 37372 42684
rect 37139 42653 37151 42656
rect 37093 42647 37151 42653
rect 37366 42644 37372 42656
rect 37424 42644 37430 42696
rect 37918 42644 37924 42696
rect 37976 42684 37982 42696
rect 38304 42693 38332 42724
rect 39850 42712 39856 42724
rect 39908 42712 39914 42764
rect 44192 42752 44220 42860
rect 44361 42755 44419 42761
rect 44361 42752 44373 42755
rect 44192 42724 44373 42752
rect 44361 42721 44373 42724
rect 44407 42752 44419 42755
rect 46566 42752 46572 42764
rect 44407 42724 46572 42752
rect 44407 42721 44419 42724
rect 44361 42715 44419 42721
rect 46566 42712 46572 42724
rect 46624 42712 46630 42764
rect 67910 42752 67916 42764
rect 67871 42724 67916 42752
rect 67910 42712 67916 42724
rect 67968 42712 67974 42764
rect 38105 42687 38163 42693
rect 38105 42684 38117 42687
rect 37976 42656 38117 42684
rect 37976 42644 37982 42656
rect 38105 42653 38117 42656
rect 38151 42653 38163 42687
rect 38105 42647 38163 42653
rect 38289 42687 38347 42693
rect 38289 42653 38301 42687
rect 38335 42653 38347 42687
rect 38289 42647 38347 42653
rect 38933 42687 38991 42693
rect 38933 42653 38945 42687
rect 38979 42653 38991 42687
rect 38933 42647 38991 42653
rect 40037 42687 40095 42693
rect 40037 42653 40049 42687
rect 40083 42684 40095 42687
rect 40126 42684 40132 42696
rect 40083 42656 40132 42684
rect 40083 42653 40095 42656
rect 40037 42647 40095 42653
rect 29914 42616 29920 42628
rect 29840 42588 29920 42616
rect 29914 42576 29920 42588
rect 29972 42616 29978 42628
rect 32401 42619 32459 42625
rect 29972 42588 32352 42616
rect 29972 42576 29978 42588
rect 23716 42520 24808 42548
rect 23716 42508 23722 42520
rect 24946 42508 24952 42560
rect 25004 42548 25010 42560
rect 25777 42551 25835 42557
rect 25777 42548 25789 42551
rect 25004 42520 25789 42548
rect 25004 42508 25010 42520
rect 25777 42517 25789 42520
rect 25823 42548 25835 42551
rect 30190 42548 30196 42560
rect 25823 42520 30196 42548
rect 25823 42517 25835 42520
rect 25777 42511 25835 42517
rect 30190 42508 30196 42520
rect 30248 42508 30254 42560
rect 31021 42551 31079 42557
rect 31021 42517 31033 42551
rect 31067 42548 31079 42551
rect 31110 42548 31116 42560
rect 31067 42520 31116 42548
rect 31067 42517 31079 42520
rect 31021 42511 31079 42517
rect 31110 42508 31116 42520
rect 31168 42508 31174 42560
rect 31754 42508 31760 42560
rect 31812 42548 31818 42560
rect 32324 42548 32352 42588
rect 32401 42585 32413 42619
rect 32447 42616 32459 42619
rect 32490 42616 32496 42628
rect 32447 42588 32496 42616
rect 32447 42585 32459 42588
rect 32401 42579 32459 42585
rect 32490 42576 32496 42588
rect 32548 42576 32554 42628
rect 33778 42616 33784 42628
rect 33739 42588 33784 42616
rect 33778 42576 33784 42588
rect 33836 42576 33842 42628
rect 34968 42619 35026 42625
rect 34968 42585 34980 42619
rect 35014 42616 35026 42619
rect 35434 42616 35440 42628
rect 35014 42588 35440 42616
rect 35014 42585 35026 42588
rect 34968 42579 35026 42585
rect 35434 42576 35440 42588
rect 35492 42576 35498 42628
rect 37642 42576 37648 42628
rect 37700 42616 37706 42628
rect 38010 42616 38016 42628
rect 37700 42588 38016 42616
rect 37700 42576 37706 42588
rect 38010 42576 38016 42588
rect 38068 42616 38074 42628
rect 38948 42616 38976 42647
rect 40126 42644 40132 42656
rect 40184 42684 40190 42696
rect 40310 42684 40316 42696
rect 40184 42656 40316 42684
rect 40184 42644 40190 42656
rect 40310 42644 40316 42656
rect 40368 42644 40374 42696
rect 41141 42687 41199 42693
rect 41141 42653 41153 42687
rect 41187 42684 41199 42687
rect 41782 42684 41788 42696
rect 41187 42656 41788 42684
rect 41187 42653 41199 42656
rect 41141 42647 41199 42653
rect 41782 42644 41788 42656
rect 41840 42644 41846 42696
rect 41874 42644 41880 42696
rect 41932 42684 41938 42696
rect 43165 42687 43223 42693
rect 43165 42684 43177 42687
rect 41932 42656 43177 42684
rect 41932 42644 41938 42656
rect 43165 42653 43177 42656
rect 43211 42653 43223 42687
rect 43165 42647 43223 42653
rect 43346 42644 43352 42696
rect 43404 42684 43410 42696
rect 45189 42687 45247 42693
rect 45189 42684 45201 42687
rect 43404 42656 45201 42684
rect 43404 42644 43410 42656
rect 45189 42653 45201 42656
rect 45235 42653 45247 42687
rect 48130 42684 48136 42696
rect 48091 42656 48136 42684
rect 45189 42647 45247 42653
rect 48130 42644 48136 42656
rect 48188 42644 48194 42696
rect 65794 42644 65800 42696
rect 65852 42684 65858 42696
rect 67269 42687 67327 42693
rect 67269 42684 67281 42687
rect 65852 42656 67281 42684
rect 65852 42644 65858 42656
rect 67269 42653 67281 42656
rect 67315 42653 67327 42687
rect 67269 42647 67327 42653
rect 38068 42588 38976 42616
rect 41408 42619 41466 42625
rect 38068 42576 38074 42588
rect 41408 42585 41420 42619
rect 41454 42616 41466 42619
rect 44082 42616 44088 42628
rect 41454 42588 43024 42616
rect 44043 42588 44088 42616
rect 41454 42585 41466 42588
rect 41408 42579 41466 42585
rect 32601 42551 32659 42557
rect 32601 42548 32613 42551
rect 31812 42520 31857 42548
rect 32324 42520 32613 42548
rect 31812 42508 31818 42520
rect 32601 42517 32613 42520
rect 32647 42548 32659 42551
rect 33962 42548 33968 42560
rect 34020 42557 34026 42560
rect 34020 42551 34039 42557
rect 32647 42520 33968 42548
rect 32647 42517 32659 42520
rect 32601 42511 32659 42517
rect 33962 42508 33968 42520
rect 34027 42517 34039 42551
rect 34020 42511 34039 42517
rect 34149 42551 34207 42557
rect 34149 42517 34161 42551
rect 34195 42548 34207 42551
rect 35710 42548 35716 42560
rect 34195 42520 35716 42548
rect 34195 42517 34207 42520
rect 34149 42511 34207 42517
rect 34020 42508 34026 42511
rect 35710 42508 35716 42520
rect 35768 42508 35774 42560
rect 36078 42548 36084 42560
rect 36039 42520 36084 42548
rect 36078 42508 36084 42520
rect 36136 42508 36142 42560
rect 37826 42508 37832 42560
rect 37884 42548 37890 42560
rect 38197 42551 38255 42557
rect 38197 42548 38209 42551
rect 37884 42520 38209 42548
rect 37884 42508 37890 42520
rect 38197 42517 38209 42520
rect 38243 42517 38255 42551
rect 38197 42511 38255 42517
rect 39758 42508 39764 42560
rect 39816 42548 39822 42560
rect 40221 42551 40279 42557
rect 40221 42548 40233 42551
rect 39816 42520 40233 42548
rect 39816 42508 39822 42520
rect 40221 42517 40233 42520
rect 40267 42517 40279 42551
rect 40221 42511 40279 42517
rect 41322 42508 41328 42560
rect 41380 42548 41386 42560
rect 42996 42557 43024 42588
rect 44082 42576 44088 42588
rect 44140 42616 44146 42628
rect 45278 42616 45284 42628
rect 44140 42588 45284 42616
rect 44140 42576 44146 42588
rect 45278 42576 45284 42588
rect 45336 42576 45342 42628
rect 42521 42551 42579 42557
rect 42521 42548 42533 42551
rect 41380 42520 42533 42548
rect 41380 42508 41386 42520
rect 42521 42517 42533 42520
rect 42567 42517 42579 42551
rect 42521 42511 42579 42517
rect 42981 42551 43039 42557
rect 42981 42517 42993 42551
rect 43027 42517 43039 42551
rect 45002 42548 45008 42560
rect 44963 42520 45008 42548
rect 42981 42511 43039 42517
rect 45002 42508 45008 42520
rect 45060 42508 45066 42560
rect 47949 42551 48007 42557
rect 47949 42517 47961 42551
rect 47995 42548 48007 42551
rect 48314 42548 48320 42560
rect 47995 42520 48320 42548
rect 47995 42517 48007 42520
rect 47949 42511 48007 42517
rect 48314 42508 48320 42520
rect 48372 42508 48378 42560
rect 1104 42458 68816 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 68816 42458
rect 1104 42384 68816 42406
rect 1946 42304 1952 42356
rect 2004 42344 2010 42356
rect 2004 42316 17448 42344
rect 2004 42304 2010 42316
rect 15004 42279 15062 42285
rect 15004 42245 15016 42279
rect 15050 42276 15062 42279
rect 15470 42276 15476 42288
rect 15050 42248 15476 42276
rect 15050 42245 15062 42248
rect 15004 42239 15062 42245
rect 15470 42236 15476 42248
rect 15528 42236 15534 42288
rect 14734 42208 14740 42220
rect 14695 42180 14740 42208
rect 14734 42168 14740 42180
rect 14792 42168 14798 42220
rect 16942 42208 16948 42220
rect 16903 42180 16948 42208
rect 16942 42168 16948 42180
rect 17000 42168 17006 42220
rect 17218 42217 17224 42220
rect 17212 42171 17224 42217
rect 17276 42208 17282 42220
rect 17420 42208 17448 42316
rect 18046 42304 18052 42356
rect 18104 42344 18110 42356
rect 18325 42347 18383 42353
rect 18325 42344 18337 42347
rect 18104 42316 18337 42344
rect 18104 42304 18110 42316
rect 18325 42313 18337 42316
rect 18371 42313 18383 42347
rect 18325 42307 18383 42313
rect 18414 42304 18420 42356
rect 18472 42344 18478 42356
rect 25038 42344 25044 42356
rect 18472 42316 25044 42344
rect 18472 42304 18478 42316
rect 25038 42304 25044 42316
rect 25096 42304 25102 42356
rect 25593 42347 25651 42353
rect 25593 42313 25605 42347
rect 25639 42344 25651 42347
rect 25866 42344 25872 42356
rect 25639 42316 25872 42344
rect 25639 42313 25651 42316
rect 25593 42307 25651 42313
rect 25866 42304 25872 42316
rect 25924 42304 25930 42356
rect 28350 42344 28356 42356
rect 28311 42316 28356 42344
rect 28350 42304 28356 42316
rect 28408 42304 28414 42356
rect 29730 42304 29736 42356
rect 29788 42344 29794 42356
rect 31018 42344 31024 42356
rect 29788 42316 31024 42344
rect 29788 42304 29794 42316
rect 31018 42304 31024 42316
rect 31076 42304 31082 42356
rect 32122 42304 32128 42356
rect 32180 42344 32186 42356
rect 34146 42344 34152 42356
rect 32180 42316 32536 42344
rect 34107 42316 34152 42344
rect 32180 42304 32186 42316
rect 17494 42236 17500 42288
rect 17552 42276 17558 42288
rect 22281 42279 22339 42285
rect 17552 42248 19748 42276
rect 17552 42236 17558 42248
rect 18782 42208 18788 42220
rect 17276 42180 17312 42208
rect 17420 42180 18000 42208
rect 18743 42180 18788 42208
rect 17218 42168 17224 42171
rect 17276 42168 17282 42180
rect 17972 42140 18000 42180
rect 18782 42168 18788 42180
rect 18840 42168 18846 42220
rect 19334 42168 19340 42220
rect 19392 42208 19398 42220
rect 19610 42208 19616 42220
rect 19392 42180 19616 42208
rect 19392 42168 19398 42180
rect 19610 42168 19616 42180
rect 19668 42168 19674 42220
rect 19720 42217 19748 42248
rect 22281 42245 22293 42279
rect 22327 42276 22339 42279
rect 30742 42276 30748 42288
rect 22327 42248 30748 42276
rect 22327 42245 22339 42248
rect 22281 42239 22339 42245
rect 30742 42236 30748 42248
rect 30800 42236 30806 42288
rect 31754 42236 31760 42288
rect 31812 42276 31818 42288
rect 32370 42279 32428 42285
rect 32370 42276 32382 42279
rect 31812 42248 32382 42276
rect 31812 42236 31818 42248
rect 32370 42245 32382 42248
rect 32416 42245 32428 42279
rect 32508 42276 32536 42316
rect 34146 42304 34152 42316
rect 34204 42304 34210 42356
rect 35434 42344 35440 42356
rect 35395 42316 35440 42344
rect 35434 42304 35440 42316
rect 35492 42304 35498 42356
rect 35526 42304 35532 42356
rect 35584 42344 35590 42356
rect 67082 42344 67088 42356
rect 35584 42316 67088 42344
rect 35584 42304 35590 42316
rect 67082 42304 67088 42316
rect 67140 42304 67146 42356
rect 34793 42279 34851 42285
rect 32508 42248 34100 42276
rect 32370 42239 32428 42245
rect 19705 42211 19763 42217
rect 19705 42177 19717 42211
rect 19751 42177 19763 42211
rect 19705 42171 19763 42177
rect 20990 42168 20996 42220
rect 21048 42208 21054 42220
rect 22649 42211 22707 42217
rect 22649 42208 22661 42211
rect 21048 42180 22661 42208
rect 21048 42168 21054 42180
rect 22649 42177 22661 42180
rect 22695 42177 22707 42211
rect 22649 42171 22707 42177
rect 23201 42211 23259 42217
rect 23201 42177 23213 42211
rect 23247 42177 23259 42211
rect 23382 42208 23388 42220
rect 23343 42180 23388 42208
rect 23201 42171 23259 42177
rect 22094 42140 22100 42152
rect 17972 42112 22100 42140
rect 22094 42100 22100 42112
rect 22152 42100 22158 42152
rect 20162 42072 20168 42084
rect 18340 42044 20168 42072
rect 16114 42004 16120 42016
rect 16075 41976 16120 42004
rect 16114 41964 16120 41976
rect 16172 42004 16178 42016
rect 18340 42004 18368 42044
rect 20162 42032 20168 42044
rect 20220 42032 20226 42084
rect 22664 42072 22692 42171
rect 23216 42140 23244 42171
rect 23382 42168 23388 42180
rect 23440 42168 23446 42220
rect 23845 42211 23903 42217
rect 23845 42177 23857 42211
rect 23891 42208 23903 42211
rect 24946 42208 24952 42220
rect 23891 42180 24716 42208
rect 24907 42180 24952 42208
rect 23891 42177 23903 42180
rect 23845 42171 23903 42177
rect 23566 42140 23572 42152
rect 23216 42112 23572 42140
rect 23566 42100 23572 42112
rect 23624 42140 23630 42152
rect 24210 42140 24216 42152
rect 23624 42112 24216 42140
rect 23624 42100 23630 42112
rect 24210 42100 24216 42112
rect 24268 42100 24274 42152
rect 24302 42072 24308 42084
rect 22664 42044 24308 42072
rect 24302 42032 24308 42044
rect 24360 42032 24366 42084
rect 24688 42072 24716 42180
rect 24946 42168 24952 42180
rect 25004 42168 25010 42220
rect 25041 42211 25099 42217
rect 25041 42177 25053 42211
rect 25087 42208 25099 42211
rect 25222 42208 25228 42220
rect 25087 42180 25228 42208
rect 25087 42177 25099 42180
rect 25041 42171 25099 42177
rect 25222 42168 25228 42180
rect 25280 42168 25286 42220
rect 25406 42168 25412 42220
rect 25464 42208 25470 42220
rect 25869 42211 25927 42217
rect 25869 42208 25881 42211
rect 25464 42180 25881 42208
rect 25464 42168 25470 42180
rect 25869 42177 25881 42180
rect 25915 42177 25927 42211
rect 26142 42208 26148 42220
rect 26103 42180 26148 42208
rect 25869 42171 25927 42177
rect 26142 42168 26148 42180
rect 26200 42168 26206 42220
rect 26970 42208 26976 42220
rect 26931 42180 26976 42208
rect 26970 42168 26976 42180
rect 27028 42168 27034 42220
rect 27433 42211 27491 42217
rect 27433 42177 27445 42211
rect 27479 42177 27491 42211
rect 27433 42171 27491 42177
rect 25958 42140 25964 42152
rect 25919 42112 25964 42140
rect 25958 42100 25964 42112
rect 26016 42100 26022 42152
rect 26329 42075 26387 42081
rect 24688 42044 26096 42072
rect 26068 42016 26096 42044
rect 26329 42041 26341 42075
rect 26375 42072 26387 42075
rect 27448 42072 27476 42171
rect 27522 42168 27528 42220
rect 27580 42208 27586 42220
rect 27801 42211 27859 42217
rect 27801 42208 27813 42211
rect 27580 42180 27813 42208
rect 27580 42168 27586 42180
rect 27801 42177 27813 42180
rect 27847 42177 27859 42211
rect 27801 42171 27859 42177
rect 28353 42211 28411 42217
rect 28353 42177 28365 42211
rect 28399 42208 28411 42211
rect 28626 42208 28632 42220
rect 28399 42180 28632 42208
rect 28399 42177 28411 42180
rect 28353 42171 28411 42177
rect 28626 42168 28632 42180
rect 28684 42168 28690 42220
rect 29086 42208 29092 42220
rect 29047 42180 29092 42208
rect 29086 42168 29092 42180
rect 29144 42168 29150 42220
rect 31110 42168 31116 42220
rect 31168 42208 31174 42220
rect 31297 42211 31355 42217
rect 31297 42208 31309 42211
rect 31168 42180 31309 42208
rect 31168 42168 31174 42180
rect 31297 42177 31309 42180
rect 31343 42208 31355 42211
rect 32766 42208 32772 42220
rect 31343 42180 32772 42208
rect 31343 42177 31355 42180
rect 31297 42171 31355 42177
rect 32766 42168 32772 42180
rect 32824 42168 32830 42220
rect 32950 42168 32956 42220
rect 33008 42208 33014 42220
rect 33962 42208 33968 42220
rect 33008 42180 33180 42208
rect 33923 42180 33968 42208
rect 33008 42168 33014 42180
rect 29178 42100 29184 42152
rect 29236 42140 29242 42152
rect 29362 42140 29368 42152
rect 29236 42112 29368 42140
rect 29236 42100 29242 42112
rect 29362 42100 29368 42112
rect 29420 42100 29426 42152
rect 31573 42143 31631 42149
rect 31573 42109 31585 42143
rect 31619 42140 31631 42143
rect 32114 42143 32172 42149
rect 32114 42140 32126 42143
rect 31619 42112 32126 42140
rect 31619 42109 31631 42112
rect 31573 42103 31631 42109
rect 32114 42109 32126 42112
rect 32160 42109 32172 42143
rect 32114 42103 32172 42109
rect 30098 42072 30104 42084
rect 26375 42044 27476 42072
rect 28184 42044 30104 42072
rect 26375 42041 26387 42044
rect 26329 42035 26387 42041
rect 16172 41976 18368 42004
rect 18969 42007 19027 42013
rect 16172 41964 16178 41976
rect 18969 41973 18981 42007
rect 19015 42004 19027 42007
rect 19242 42004 19248 42016
rect 19015 41976 19248 42004
rect 19015 41973 19027 41976
rect 18969 41967 19027 41973
rect 19242 41964 19248 41976
rect 19300 41964 19306 42016
rect 19889 42007 19947 42013
rect 19889 41973 19901 42007
rect 19935 42004 19947 42007
rect 19978 42004 19984 42016
rect 19935 41976 19984 42004
rect 19935 41973 19947 41976
rect 19889 41967 19947 41973
rect 19978 41964 19984 41976
rect 20036 41964 20042 42016
rect 24026 42004 24032 42016
rect 23987 41976 24032 42004
rect 24026 41964 24032 41976
rect 24084 41964 24090 42016
rect 24578 41964 24584 42016
rect 24636 42004 24642 42016
rect 25225 42007 25283 42013
rect 25225 42004 25237 42007
rect 24636 41976 25237 42004
rect 24636 41964 24642 41976
rect 25225 41973 25237 41976
rect 25271 41973 25283 42007
rect 25866 42004 25872 42016
rect 25827 41976 25872 42004
rect 25225 41967 25283 41973
rect 25866 41964 25872 41976
rect 25924 41964 25930 42016
rect 26050 41964 26056 42016
rect 26108 42004 26114 42016
rect 28184 42004 28212 42044
rect 30098 42032 30104 42044
rect 30156 42032 30162 42084
rect 33152 42072 33180 42180
rect 33962 42168 33968 42180
rect 34020 42168 34026 42220
rect 34072 42208 34100 42248
rect 34793 42245 34805 42279
rect 34839 42276 34851 42279
rect 37918 42276 37924 42288
rect 34839 42248 37924 42276
rect 34839 42245 34851 42248
rect 34793 42239 34851 42245
rect 37918 42236 37924 42248
rect 37976 42236 37982 42288
rect 41601 42279 41659 42285
rect 41601 42245 41613 42279
rect 41647 42276 41659 42279
rect 41874 42276 41880 42288
rect 41647 42248 41880 42276
rect 41647 42245 41659 42248
rect 41601 42239 41659 42245
rect 41874 42236 41880 42248
rect 41932 42236 41938 42288
rect 43346 42276 43352 42288
rect 43307 42248 43352 42276
rect 43346 42236 43352 42248
rect 43404 42236 43410 42288
rect 44076 42279 44134 42285
rect 44076 42245 44088 42279
rect 44122 42276 44134 42279
rect 45002 42276 45008 42288
rect 44122 42248 45008 42276
rect 44122 42245 44134 42248
rect 44076 42239 44134 42245
rect 45002 42236 45008 42248
rect 45060 42236 45066 42288
rect 35526 42208 35532 42220
rect 34072 42180 35532 42208
rect 35526 42168 35532 42180
rect 35584 42168 35590 42220
rect 35621 42211 35679 42217
rect 35621 42177 35633 42211
rect 35667 42208 35679 42211
rect 35710 42208 35716 42220
rect 35667 42180 35716 42208
rect 35667 42177 35679 42180
rect 35621 42171 35679 42177
rect 35710 42168 35716 42180
rect 35768 42168 35774 42220
rect 35986 42168 35992 42220
rect 36044 42208 36050 42220
rect 36357 42211 36415 42217
rect 36357 42208 36369 42211
rect 36044 42180 36369 42208
rect 36044 42168 36050 42180
rect 36357 42177 36369 42180
rect 36403 42177 36415 42211
rect 36538 42208 36544 42220
rect 36499 42180 36544 42208
rect 36357 42171 36415 42177
rect 36538 42168 36544 42180
rect 36596 42168 36602 42220
rect 37277 42211 37335 42217
rect 37277 42177 37289 42211
rect 37323 42177 37335 42211
rect 37277 42171 37335 42177
rect 33410 42100 33416 42152
rect 33468 42140 33474 42152
rect 33778 42140 33784 42152
rect 33468 42112 33784 42140
rect 33468 42100 33474 42112
rect 33778 42100 33784 42112
rect 33836 42140 33842 42152
rect 36078 42140 36084 42152
rect 33836 42112 36084 42140
rect 33836 42100 33842 42112
rect 36078 42100 36084 42112
rect 36136 42100 36142 42152
rect 37292 42140 37320 42171
rect 37366 42168 37372 42220
rect 37424 42208 37430 42220
rect 37461 42211 37519 42217
rect 37461 42208 37473 42211
rect 37424 42180 37473 42208
rect 37424 42168 37430 42180
rect 37461 42177 37473 42180
rect 37507 42177 37519 42211
rect 37461 42171 37519 42177
rect 38565 42211 38623 42217
rect 38565 42177 38577 42211
rect 38611 42208 38623 42211
rect 39574 42208 39580 42220
rect 38611 42180 39580 42208
rect 38611 42177 38623 42180
rect 38565 42171 38623 42177
rect 39574 42168 39580 42180
rect 39632 42168 39638 42220
rect 39758 42208 39764 42220
rect 39719 42180 39764 42208
rect 39758 42168 39764 42180
rect 39816 42168 39822 42220
rect 41322 42208 41328 42220
rect 41283 42180 41328 42208
rect 41322 42168 41328 42180
rect 41380 42168 41386 42220
rect 41417 42211 41475 42217
rect 41417 42177 41429 42211
rect 41463 42208 41475 42211
rect 41690 42208 41696 42220
rect 41463 42180 41696 42208
rect 41463 42177 41475 42180
rect 41417 42171 41475 42177
rect 41690 42168 41696 42180
rect 41748 42208 41754 42220
rect 43165 42211 43223 42217
rect 43165 42208 43177 42211
rect 41748 42180 43177 42208
rect 41748 42168 41754 42180
rect 43165 42177 43177 42180
rect 43211 42208 43223 42211
rect 43622 42208 43628 42220
rect 43211 42180 43628 42208
rect 43211 42177 43223 42180
rect 43165 42171 43223 42177
rect 43622 42168 43628 42180
rect 43680 42168 43686 42220
rect 43806 42208 43812 42220
rect 43767 42180 43812 42208
rect 43806 42168 43812 42180
rect 43864 42168 43870 42220
rect 65794 42208 65800 42220
rect 65755 42180 65800 42208
rect 65794 42168 65800 42180
rect 65852 42168 65858 42220
rect 36188 42112 37320 42140
rect 38657 42143 38715 42149
rect 36188 42072 36216 42112
rect 38657 42109 38669 42143
rect 38703 42109 38715 42143
rect 38657 42103 38715 42109
rect 38749 42143 38807 42149
rect 38749 42109 38761 42143
rect 38795 42109 38807 42143
rect 38749 42103 38807 42109
rect 38841 42143 38899 42149
rect 38841 42109 38853 42143
rect 38887 42140 38899 42143
rect 39022 42140 39028 42152
rect 38887 42112 39028 42140
rect 38887 42109 38899 42112
rect 38841 42103 38899 42109
rect 33152 42044 36216 42072
rect 36725 42075 36783 42081
rect 36725 42041 36737 42075
rect 36771 42072 36783 42075
rect 38672 42072 38700 42103
rect 36771 42044 38700 42072
rect 38764 42072 38792 42103
rect 39022 42100 39028 42112
rect 39080 42140 39086 42152
rect 42426 42140 42432 42152
rect 39080 42112 42432 42140
rect 39080 42100 39086 42112
rect 42426 42100 42432 42112
rect 42484 42100 42490 42152
rect 42981 42143 43039 42149
rect 42981 42109 42993 42143
rect 43027 42140 43039 42143
rect 48590 42140 48596 42152
rect 43027 42112 43852 42140
rect 48551 42112 48596 42140
rect 43027 42109 43039 42112
rect 42981 42103 43039 42109
rect 43180 42084 43208 42112
rect 38930 42072 38936 42084
rect 38764 42044 38936 42072
rect 36771 42041 36783 42044
rect 36725 42035 36783 42041
rect 38930 42032 38936 42044
rect 38988 42072 38994 42084
rect 39206 42072 39212 42084
rect 38988 42044 39212 42072
rect 38988 42032 38994 42044
rect 39206 42032 39212 42044
rect 39264 42032 39270 42084
rect 39390 42032 39396 42084
rect 39448 42072 39454 42084
rect 39577 42075 39635 42081
rect 39577 42072 39589 42075
rect 39448 42044 39589 42072
rect 39448 42032 39454 42044
rect 39577 42041 39589 42044
rect 39623 42041 39635 42075
rect 39577 42035 39635 42041
rect 43162 42032 43168 42084
rect 43220 42032 43226 42084
rect 28902 42004 28908 42016
rect 26108 41976 28212 42004
rect 28863 41976 28908 42004
rect 26108 41964 26114 41976
rect 28902 41964 28908 41976
rect 28960 41964 28966 42016
rect 29178 41964 29184 42016
rect 29236 42004 29242 42016
rect 32122 42004 32128 42016
rect 29236 41976 32128 42004
rect 29236 41964 29242 41976
rect 32122 41964 32128 41976
rect 32180 41964 32186 42016
rect 32490 41964 32496 42016
rect 32548 42004 32554 42016
rect 33505 42007 33563 42013
rect 33505 42004 33517 42007
rect 32548 41976 33517 42004
rect 32548 41964 32554 41976
rect 33505 41973 33517 41976
rect 33551 41973 33563 42007
rect 33505 41967 33563 41973
rect 34790 41964 34796 42016
rect 34848 42004 34854 42016
rect 34885 42007 34943 42013
rect 34885 42004 34897 42007
rect 34848 41976 34897 42004
rect 34848 41964 34854 41976
rect 34885 41973 34897 41976
rect 34931 41973 34943 42007
rect 37642 42004 37648 42016
rect 37603 41976 37648 42004
rect 34885 41967 34943 41973
rect 37642 41964 37648 41976
rect 37700 41964 37706 42016
rect 38381 42007 38439 42013
rect 38381 41973 38393 42007
rect 38427 42004 38439 42007
rect 38838 42004 38844 42016
rect 38427 41976 38844 42004
rect 38427 41973 38439 41976
rect 38381 41967 38439 41973
rect 38838 41964 38844 41976
rect 38896 41964 38902 42016
rect 43824 42004 43852 42112
rect 48590 42100 48596 42112
rect 48648 42100 48654 42152
rect 48777 42143 48835 42149
rect 48777 42109 48789 42143
rect 48823 42140 48835 42143
rect 49418 42140 49424 42152
rect 48823 42112 49424 42140
rect 48823 42109 48835 42112
rect 48777 42103 48835 42109
rect 49418 42100 49424 42112
rect 49476 42100 49482 42152
rect 50433 42143 50491 42149
rect 50433 42109 50445 42143
rect 50479 42140 50491 42143
rect 64874 42140 64880 42152
rect 50479 42112 64880 42140
rect 50479 42109 50491 42112
rect 50433 42103 50491 42109
rect 64874 42100 64880 42112
rect 64932 42100 64938 42152
rect 65978 42140 65984 42152
rect 65939 42112 65984 42140
rect 65978 42100 65984 42112
rect 66036 42100 66042 42152
rect 67542 42140 67548 42152
rect 67503 42112 67548 42140
rect 67542 42100 67548 42112
rect 67600 42100 67606 42152
rect 45189 42007 45247 42013
rect 45189 42004 45201 42007
rect 43824 41976 45201 42004
rect 45189 41973 45201 41976
rect 45235 41973 45247 42007
rect 45189 41967 45247 41973
rect 1104 41914 68816 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 65654 41914
rect 65706 41862 65718 41914
rect 65770 41862 65782 41914
rect 65834 41862 65846 41914
rect 65898 41862 65910 41914
rect 65962 41862 68816 41914
rect 1104 41840 68816 41862
rect 15746 41800 15752 41812
rect 15707 41772 15752 41800
rect 15746 41760 15752 41772
rect 15804 41760 15810 41812
rect 17037 41803 17095 41809
rect 17037 41769 17049 41803
rect 17083 41800 17095 41803
rect 17589 41803 17647 41809
rect 17589 41800 17601 41803
rect 17083 41772 17601 41800
rect 17083 41769 17095 41772
rect 17037 41763 17095 41769
rect 17589 41769 17601 41772
rect 17635 41800 17647 41803
rect 17635 41772 19104 41800
rect 17635 41769 17647 41772
rect 17589 41763 17647 41769
rect 14826 41692 14832 41744
rect 14884 41732 14890 41744
rect 17773 41735 17831 41741
rect 14884 41704 16574 41732
rect 14884 41692 14890 41704
rect 15381 41667 15439 41673
rect 15381 41633 15393 41667
rect 15427 41664 15439 41667
rect 16114 41664 16120 41676
rect 15427 41636 16120 41664
rect 15427 41633 15439 41636
rect 15381 41627 15439 41633
rect 16114 41624 16120 41636
rect 16172 41624 16178 41676
rect 16546 41664 16574 41704
rect 17773 41701 17785 41735
rect 17819 41732 17831 41735
rect 18414 41732 18420 41744
rect 17819 41704 18420 41732
rect 17819 41701 17831 41704
rect 17773 41695 17831 41701
rect 18414 41692 18420 41704
rect 18472 41692 18478 41744
rect 17405 41667 17463 41673
rect 17405 41664 17417 41667
rect 16546 41636 17417 41664
rect 17405 41633 17417 41636
rect 17451 41633 17463 41667
rect 17405 41627 17463 41633
rect 15562 41596 15568 41608
rect 15523 41568 15568 41596
rect 15562 41556 15568 41568
rect 15620 41556 15626 41608
rect 17586 41596 17592 41608
rect 17547 41568 17592 41596
rect 17586 41556 17592 41568
rect 17644 41556 17650 41608
rect 19076 41596 19104 41772
rect 19610 41760 19616 41812
rect 19668 41800 19674 41812
rect 20625 41803 20683 41809
rect 20625 41800 20637 41803
rect 19668 41772 20637 41800
rect 19668 41760 19674 41772
rect 20625 41769 20637 41772
rect 20671 41769 20683 41803
rect 23569 41803 23627 41809
rect 20625 41763 20683 41769
rect 20732 41772 22048 41800
rect 19242 41664 19248 41676
rect 19203 41636 19248 41664
rect 19242 41624 19248 41636
rect 19300 41624 19306 41676
rect 20732 41596 20760 41772
rect 22020 41732 22048 41772
rect 23569 41769 23581 41803
rect 23615 41800 23627 41803
rect 23658 41800 23664 41812
rect 23615 41772 23664 41800
rect 23615 41769 23627 41772
rect 23569 41763 23627 41769
rect 23658 41760 23664 41772
rect 23716 41760 23722 41812
rect 24397 41803 24455 41809
rect 24397 41769 24409 41803
rect 24443 41800 24455 41803
rect 24486 41800 24492 41812
rect 24443 41772 24492 41800
rect 24443 41769 24455 41772
rect 24397 41763 24455 41769
rect 24486 41760 24492 41772
rect 24544 41760 24550 41812
rect 25774 41800 25780 41812
rect 25735 41772 25780 41800
rect 25774 41760 25780 41772
rect 25832 41800 25838 41812
rect 26326 41800 26332 41812
rect 25832 41772 26332 41800
rect 25832 41760 25838 41772
rect 26326 41760 26332 41772
rect 26384 41760 26390 41812
rect 26421 41803 26479 41809
rect 26421 41769 26433 41803
rect 26467 41800 26479 41803
rect 26510 41800 26516 41812
rect 26467 41772 26516 41800
rect 26467 41769 26479 41772
rect 26421 41763 26479 41769
rect 26510 41760 26516 41772
rect 26568 41760 26574 41812
rect 26605 41803 26663 41809
rect 26605 41769 26617 41803
rect 26651 41800 26663 41803
rect 27522 41800 27528 41812
rect 26651 41772 27528 41800
rect 26651 41769 26663 41772
rect 26605 41763 26663 41769
rect 27522 41760 27528 41772
rect 27580 41760 27586 41812
rect 58710 41800 58716 41812
rect 27632 41772 58716 41800
rect 27632 41732 27660 41772
rect 58710 41760 58716 41772
rect 58768 41760 58774 41812
rect 65978 41760 65984 41812
rect 66036 41800 66042 41812
rect 67637 41803 67695 41809
rect 67637 41800 67649 41803
rect 66036 41772 67649 41800
rect 66036 41760 66042 41772
rect 67637 41769 67649 41772
rect 67683 41769 67695 41803
rect 67637 41763 67695 41769
rect 28994 41732 29000 41744
rect 22020 41704 27660 41732
rect 28907 41704 29000 41732
rect 28994 41692 29000 41704
rect 29052 41732 29058 41744
rect 29454 41732 29460 41744
rect 29052 41704 29460 41732
rect 29052 41692 29058 41704
rect 29454 41692 29460 41704
rect 29512 41692 29518 41744
rect 31018 41692 31024 41744
rect 31076 41732 31082 41744
rect 37274 41732 37280 41744
rect 31076 41704 37280 41732
rect 31076 41692 31082 41704
rect 37274 41692 37280 41704
rect 37332 41692 37338 41744
rect 39022 41692 39028 41744
rect 39080 41732 39086 41744
rect 46290 41732 46296 41744
rect 39080 41704 46296 41732
rect 39080 41692 39086 41704
rect 22094 41624 22100 41676
rect 22152 41664 22158 41676
rect 26237 41667 26295 41673
rect 26237 41664 26249 41667
rect 22152 41636 26249 41664
rect 22152 41624 22158 41636
rect 26237 41633 26249 41636
rect 26283 41633 26295 41667
rect 32309 41667 32367 41673
rect 32309 41664 32321 41667
rect 26237 41627 26295 41633
rect 31726 41636 32321 41664
rect 19076 41568 20760 41596
rect 21085 41599 21143 41605
rect 21085 41565 21097 41599
rect 21131 41596 21143 41599
rect 21174 41596 21180 41608
rect 21131 41568 21180 41596
rect 21131 41565 21143 41568
rect 21085 41559 21143 41565
rect 21174 41556 21180 41568
rect 21232 41556 21238 41608
rect 23385 41599 23443 41605
rect 23385 41565 23397 41599
rect 23431 41596 23443 41599
rect 23566 41596 23572 41608
rect 23431 41568 23572 41596
rect 23431 41565 23443 41568
rect 23385 41559 23443 41565
rect 23566 41556 23572 41568
rect 23624 41556 23630 41608
rect 24578 41596 24584 41608
rect 24539 41568 24584 41596
rect 24578 41556 24584 41568
rect 24636 41556 24642 41608
rect 26145 41599 26203 41605
rect 26145 41565 26157 41599
rect 26191 41596 26203 41599
rect 26191 41568 26280 41596
rect 26191 41565 26203 41568
rect 26145 41559 26203 41565
rect 17313 41531 17371 41537
rect 17313 41497 17325 41531
rect 17359 41528 17371 41531
rect 17678 41528 17684 41540
rect 17359 41500 17684 41528
rect 17359 41497 17371 41500
rect 17313 41491 17371 41497
rect 17678 41488 17684 41500
rect 17736 41488 17742 41540
rect 19512 41531 19570 41537
rect 19512 41497 19524 41531
rect 19558 41497 19570 41531
rect 19512 41491 19570 41497
rect 21352 41531 21410 41537
rect 21352 41497 21364 41531
rect 21398 41528 21410 41531
rect 21818 41528 21824 41540
rect 21398 41500 21824 41528
rect 21398 41497 21410 41500
rect 21352 41491 21410 41497
rect 19426 41420 19432 41472
rect 19484 41460 19490 41472
rect 19536 41460 19564 41491
rect 21818 41488 21824 41500
rect 21876 41488 21882 41540
rect 19484 41432 19564 41460
rect 19484 41420 19490 41432
rect 21910 41420 21916 41472
rect 21968 41460 21974 41472
rect 22465 41463 22523 41469
rect 22465 41460 22477 41463
rect 21968 41432 22477 41460
rect 21968 41420 21974 41432
rect 22465 41429 22477 41432
rect 22511 41429 22523 41463
rect 22465 41423 22523 41429
rect 23106 41420 23112 41472
rect 23164 41460 23170 41472
rect 23382 41460 23388 41472
rect 23164 41432 23388 41460
rect 23164 41420 23170 41432
rect 23382 41420 23388 41432
rect 23440 41420 23446 41472
rect 26252 41460 26280 41568
rect 26326 41556 26332 41608
rect 26384 41596 26390 41608
rect 26421 41599 26479 41605
rect 26421 41596 26433 41599
rect 26384 41568 26433 41596
rect 26384 41556 26390 41568
rect 26421 41565 26433 41568
rect 26467 41565 26479 41599
rect 26421 41559 26479 41565
rect 27617 41599 27675 41605
rect 27617 41565 27629 41599
rect 27663 41596 27675 41599
rect 27706 41596 27712 41608
rect 27663 41568 27712 41596
rect 27663 41565 27675 41568
rect 27617 41559 27675 41565
rect 27706 41556 27712 41568
rect 27764 41556 27770 41608
rect 28166 41556 28172 41608
rect 28224 41596 28230 41608
rect 28224 41568 29868 41596
rect 28224 41556 28230 41568
rect 27884 41531 27942 41537
rect 27884 41497 27896 41531
rect 27930 41528 27942 41531
rect 28902 41528 28908 41540
rect 27930 41500 28908 41528
rect 27930 41497 27942 41500
rect 27884 41491 27942 41497
rect 28902 41488 28908 41500
rect 28960 41488 28966 41540
rect 29840 41528 29868 41568
rect 29914 41556 29920 41608
rect 29972 41596 29978 41608
rect 31726 41596 31754 41636
rect 32309 41633 32321 41636
rect 32355 41664 32367 41667
rect 38378 41664 38384 41676
rect 32355 41636 38384 41664
rect 32355 41633 32367 41636
rect 32309 41627 32367 41633
rect 38378 41624 38384 41636
rect 38436 41624 38442 41676
rect 39040 41664 39068 41692
rect 39040 41636 39151 41664
rect 29972 41568 30017 41596
rect 30116 41568 31754 41596
rect 29972 41556 29978 41568
rect 30116 41528 30144 41568
rect 32766 41556 32772 41608
rect 32824 41596 32830 41608
rect 33229 41599 33287 41605
rect 33229 41596 33241 41599
rect 32824 41568 33241 41596
rect 32824 41556 32830 41568
rect 33229 41565 33241 41568
rect 33275 41596 33287 41599
rect 33962 41596 33968 41608
rect 33275 41568 33968 41596
rect 33275 41565 33287 41568
rect 33229 41559 33287 41565
rect 33962 41556 33968 41568
rect 34020 41556 34026 41608
rect 35434 41596 35440 41608
rect 35395 41568 35440 41596
rect 35434 41556 35440 41568
rect 35492 41556 35498 41608
rect 35526 41556 35532 41608
rect 35584 41596 35590 41608
rect 37185 41599 37243 41605
rect 37185 41596 37197 41599
rect 35584 41568 37197 41596
rect 35584 41556 35590 41568
rect 37185 41565 37197 41568
rect 37231 41565 37243 41599
rect 37185 41559 37243 41565
rect 37553 41599 37611 41605
rect 37553 41565 37565 41599
rect 37599 41596 37611 41599
rect 38286 41596 38292 41608
rect 37599 41568 38292 41596
rect 37599 41565 37611 41568
rect 37553 41559 37611 41565
rect 38286 41556 38292 41568
rect 38344 41556 38350 41608
rect 38654 41605 38660 41608
rect 38611 41599 38660 41605
rect 38611 41565 38623 41599
rect 38657 41565 38660 41599
rect 38611 41559 38660 41565
rect 38654 41556 38660 41559
rect 38712 41556 38718 41608
rect 38749 41599 38807 41605
rect 38749 41565 38761 41599
rect 38795 41565 38807 41599
rect 38749 41559 38807 41565
rect 29840 41500 30144 41528
rect 30184 41531 30242 41537
rect 30184 41497 30196 41531
rect 30230 41528 30242 41531
rect 30650 41528 30656 41540
rect 30230 41500 30656 41528
rect 30230 41497 30242 41500
rect 30184 41491 30242 41497
rect 30650 41488 30656 41500
rect 30708 41488 30714 41540
rect 32125 41531 32183 41537
rect 32125 41497 32137 41531
rect 32171 41528 32183 41531
rect 34790 41528 34796 41540
rect 32171 41500 34796 41528
rect 32171 41497 32183 41500
rect 32125 41491 32183 41497
rect 34790 41488 34796 41500
rect 34848 41488 34854 41540
rect 36538 41528 36544 41540
rect 36451 41500 36544 41528
rect 36538 41488 36544 41500
rect 36596 41528 36602 41540
rect 37274 41528 37280 41540
rect 36596 41500 37280 41528
rect 36596 41488 36602 41500
rect 37274 41488 37280 41500
rect 37332 41488 37338 41540
rect 37369 41531 37427 41537
rect 37369 41497 37381 41531
rect 37415 41528 37427 41531
rect 38102 41528 38108 41540
rect 37415 41500 38108 41528
rect 37415 41497 37427 41500
rect 37369 41491 37427 41497
rect 38102 41488 38108 41500
rect 38160 41488 38166 41540
rect 38764 41528 38792 41559
rect 38838 41556 38844 41608
rect 38896 41605 38902 41608
rect 38896 41596 38904 41605
rect 39025 41599 39083 41605
rect 38896 41568 38941 41596
rect 38896 41559 38904 41568
rect 39025 41565 39037 41599
rect 39071 41593 39083 41599
rect 39123 41593 39151 41636
rect 39574 41624 39580 41676
rect 39632 41664 39638 41676
rect 42242 41673 42248 41676
rect 41417 41667 41475 41673
rect 41417 41664 41429 41667
rect 39632 41636 41429 41664
rect 39632 41624 39638 41636
rect 41417 41633 41429 41636
rect 41463 41633 41475 41667
rect 41417 41627 41475 41633
rect 42234 41667 42248 41673
rect 42234 41633 42246 41667
rect 42300 41664 42306 41676
rect 42300 41636 42334 41664
rect 42234 41627 42248 41633
rect 42242 41624 42248 41627
rect 42300 41624 42306 41636
rect 42426 41624 42432 41676
rect 42484 41664 42490 41676
rect 43349 41667 43407 41673
rect 43349 41664 43361 41667
rect 42484 41636 42529 41664
rect 42904 41636 43361 41664
rect 42484 41624 42490 41636
rect 39071 41565 39151 41593
rect 41233 41599 41291 41605
rect 41233 41565 41245 41599
rect 41279 41596 41291 41599
rect 41322 41596 41328 41608
rect 41279 41568 41328 41596
rect 41279 41565 41291 41568
rect 39025 41559 39083 41565
rect 41233 41559 41291 41565
rect 38896 41556 38902 41559
rect 41322 41556 41328 41568
rect 41380 41556 41386 41608
rect 42153 41599 42211 41605
rect 42153 41565 42165 41599
rect 42199 41565 42211 41599
rect 42334 41596 42340 41608
rect 42295 41568 42340 41596
rect 42153 41559 42211 41565
rect 38930 41528 38936 41540
rect 38764 41500 38936 41528
rect 38930 41488 38936 41500
rect 38988 41488 38994 41540
rect 41049 41531 41107 41537
rect 41049 41497 41061 41531
rect 41095 41497 41107 41531
rect 41049 41491 41107 41497
rect 26973 41463 27031 41469
rect 26973 41460 26985 41463
rect 26252 41432 26985 41460
rect 26973 41429 26985 41432
rect 27019 41460 27031 41463
rect 29178 41460 29184 41472
rect 27019 41432 29184 41460
rect 27019 41429 27031 41432
rect 26973 41423 27031 41429
rect 29178 41420 29184 41432
rect 29236 41420 29242 41472
rect 31294 41460 31300 41472
rect 31255 41432 31300 41460
rect 31294 41420 31300 41432
rect 31352 41420 31358 41472
rect 32766 41420 32772 41472
rect 32824 41460 32830 41472
rect 33321 41463 33379 41469
rect 33321 41460 33333 41463
rect 32824 41432 33333 41460
rect 32824 41420 32830 41432
rect 33321 41429 33333 41432
rect 33367 41429 33379 41463
rect 35250 41460 35256 41472
rect 35211 41432 35256 41460
rect 33321 41423 33379 41429
rect 35250 41420 35256 41432
rect 35308 41420 35314 41472
rect 36633 41463 36691 41469
rect 36633 41429 36645 41463
rect 36679 41460 36691 41463
rect 37458 41460 37464 41472
rect 36679 41432 37464 41460
rect 36679 41429 36691 41432
rect 36633 41423 36691 41429
rect 37458 41420 37464 41432
rect 37516 41460 37522 41472
rect 37734 41460 37740 41472
rect 37516 41432 37740 41460
rect 37516 41420 37522 41432
rect 37734 41420 37740 41432
rect 37792 41420 37798 41472
rect 38381 41463 38439 41469
rect 38381 41429 38393 41463
rect 38427 41460 38439 41463
rect 39022 41460 39028 41472
rect 38427 41432 39028 41460
rect 38427 41429 38439 41432
rect 38381 41423 38439 41429
rect 39022 41420 39028 41432
rect 39080 41420 39086 41472
rect 41064 41460 41092 41491
rect 41506 41488 41512 41540
rect 41564 41488 41570 41540
rect 42168 41528 42196 41559
rect 42334 41556 42340 41568
rect 42392 41556 42398 41608
rect 42904 41596 42932 41636
rect 43349 41633 43361 41636
rect 43395 41633 43407 41667
rect 43349 41627 43407 41633
rect 45370 41624 45376 41676
rect 45428 41664 45434 41676
rect 45428 41636 45600 41664
rect 45428 41624 45434 41636
rect 43162 41596 43168 41608
rect 42536 41568 42932 41596
rect 43123 41568 43168 41596
rect 42536 41528 42564 41568
rect 43162 41556 43168 41568
rect 43220 41556 43226 41608
rect 45462 41596 45468 41608
rect 45423 41568 45468 41596
rect 45462 41556 45468 41568
rect 45520 41556 45526 41608
rect 45572 41605 45600 41636
rect 45557 41599 45615 41605
rect 45557 41565 45569 41599
rect 45603 41565 45615 41599
rect 45557 41559 45615 41565
rect 45649 41599 45707 41605
rect 45649 41565 45661 41599
rect 45695 41596 45707 41599
rect 45738 41596 45744 41608
rect 45695 41568 45744 41596
rect 45695 41565 45707 41568
rect 45649 41559 45707 41565
rect 45738 41556 45744 41568
rect 45796 41556 45802 41608
rect 45848 41605 45876 41704
rect 46290 41692 46296 41704
rect 46348 41692 46354 41744
rect 49418 41732 49424 41744
rect 49379 41704 49424 41732
rect 49418 41692 49424 41704
rect 49476 41692 49482 41744
rect 45833 41599 45891 41605
rect 45833 41565 45845 41599
rect 45879 41565 45891 41599
rect 45833 41559 45891 41565
rect 46293 41599 46351 41605
rect 46293 41565 46305 41599
rect 46339 41596 46351 41599
rect 48685 41599 48743 41605
rect 46339 41568 46704 41596
rect 46339 41565 46351 41568
rect 46293 41559 46351 41565
rect 46676 41540 46704 41568
rect 48685 41565 48697 41599
rect 48731 41596 48743 41599
rect 48774 41596 48780 41608
rect 48731 41568 48780 41596
rect 48731 41565 48743 41568
rect 48685 41559 48743 41565
rect 48774 41556 48780 41568
rect 48832 41596 48838 41608
rect 49329 41599 49387 41605
rect 49329 41596 49341 41599
rect 48832 41568 49341 41596
rect 48832 41556 48838 41568
rect 49329 41565 49341 41568
rect 49375 41565 49387 41599
rect 49329 41559 49387 41565
rect 66990 41556 66996 41608
rect 67048 41596 67054 41608
rect 67545 41599 67603 41605
rect 67545 41596 67557 41599
rect 67048 41568 67557 41596
rect 67048 41556 67054 41568
rect 67545 41565 67557 41568
rect 67591 41565 67603 41599
rect 67545 41559 67603 41565
rect 42168 41500 42564 41528
rect 42886 41488 42892 41540
rect 42944 41528 42950 41540
rect 42981 41531 43039 41537
rect 42981 41528 42993 41531
rect 42944 41500 42993 41528
rect 42944 41488 42950 41500
rect 42981 41497 42993 41500
rect 43027 41497 43039 41531
rect 46538 41531 46596 41537
rect 46538 41528 46550 41531
rect 42981 41491 43039 41497
rect 45572 41500 46550 41528
rect 41524 41460 41552 41488
rect 41966 41460 41972 41472
rect 41064 41432 41552 41460
rect 41927 41432 41972 41460
rect 41966 41420 41972 41432
rect 42024 41420 42030 41472
rect 42334 41420 42340 41472
rect 42392 41460 42398 41472
rect 42794 41460 42800 41472
rect 42392 41432 42800 41460
rect 42392 41420 42398 41432
rect 42794 41420 42800 41432
rect 42852 41420 42858 41472
rect 45189 41463 45247 41469
rect 45189 41429 45201 41463
rect 45235 41460 45247 41463
rect 45572 41460 45600 41500
rect 46538 41497 46550 41500
rect 46584 41497 46596 41531
rect 46538 41491 46596 41497
rect 46658 41488 46664 41540
rect 46716 41488 46722 41540
rect 45235 41432 45600 41460
rect 45235 41429 45247 41432
rect 45189 41423 45247 41429
rect 45646 41420 45652 41472
rect 45704 41460 45710 41472
rect 47673 41463 47731 41469
rect 47673 41460 47685 41463
rect 45704 41432 47685 41460
rect 45704 41420 45710 41432
rect 47673 41429 47685 41432
rect 47719 41460 47731 41463
rect 48590 41460 48596 41472
rect 47719 41432 48596 41460
rect 47719 41429 47731 41432
rect 47673 41423 47731 41429
rect 48590 41420 48596 41432
rect 48648 41420 48654 41472
rect 48777 41463 48835 41469
rect 48777 41429 48789 41463
rect 48823 41460 48835 41463
rect 48866 41460 48872 41472
rect 48823 41432 48872 41460
rect 48823 41429 48835 41432
rect 48777 41423 48835 41429
rect 48866 41420 48872 41432
rect 48924 41420 48930 41472
rect 1104 41370 68816 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 68816 41370
rect 1104 41296 68816 41318
rect 17218 41216 17224 41268
rect 17276 41256 17282 41268
rect 17405 41259 17463 41265
rect 17405 41256 17417 41259
rect 17276 41228 17417 41256
rect 17276 41216 17282 41228
rect 17405 41225 17417 41228
rect 17451 41225 17463 41259
rect 19426 41256 19432 41268
rect 19387 41228 19432 41256
rect 17405 41219 17463 41225
rect 19426 41216 19432 41228
rect 19484 41216 19490 41268
rect 21818 41256 21824 41268
rect 21779 41228 21824 41256
rect 21818 41216 21824 41228
rect 21876 41216 21882 41268
rect 23290 41216 23296 41268
rect 23348 41256 23354 41268
rect 23661 41259 23719 41265
rect 23661 41256 23673 41259
rect 23348 41228 23673 41256
rect 23348 41216 23354 41228
rect 23661 41225 23673 41228
rect 23707 41256 23719 41259
rect 28721 41259 28779 41265
rect 23707 41228 28672 41256
rect 23707 41225 23719 41228
rect 23661 41219 23719 41225
rect 23385 41191 23443 41197
rect 23385 41157 23397 41191
rect 23431 41188 23443 41191
rect 23474 41188 23480 41200
rect 23431 41160 23480 41188
rect 23431 41157 23443 41160
rect 23385 41151 23443 41157
rect 23474 41148 23480 41160
rect 23532 41148 23538 41200
rect 24026 41148 24032 41200
rect 24084 41188 24090 41200
rect 27706 41188 27712 41200
rect 24084 41160 25452 41188
rect 27667 41160 27712 41188
rect 24084 41148 24090 41160
rect 17589 41123 17647 41129
rect 17589 41089 17601 41123
rect 17635 41120 17647 41123
rect 17954 41120 17960 41132
rect 17635 41092 17960 41120
rect 17635 41089 17647 41092
rect 17589 41083 17647 41089
rect 17954 41080 17960 41092
rect 18012 41080 18018 41132
rect 19613 41123 19671 41129
rect 19613 41089 19625 41123
rect 19659 41120 19671 41123
rect 19978 41120 19984 41132
rect 19659 41092 19984 41120
rect 19659 41089 19671 41092
rect 19613 41083 19671 41089
rect 19978 41080 19984 41092
rect 20036 41080 20042 41132
rect 22097 41123 22155 41129
rect 22097 41089 22109 41123
rect 22143 41089 22155 41123
rect 22189 41123 22247 41129
rect 22189 41116 22201 41123
rect 22235 41116 22247 41123
rect 22097 41083 22155 41089
rect 19242 41012 19248 41064
rect 19300 41052 19306 41064
rect 21910 41052 21916 41064
rect 19300 41024 21916 41052
rect 19300 41012 19306 41024
rect 21910 41012 21916 41024
rect 21968 41012 21974 41064
rect 21928 40984 21956 41012
rect 22112 40984 22140 41083
rect 22186 41064 22192 41116
rect 22244 41064 22250 41116
rect 22278 41080 22284 41132
rect 22336 41120 22342 41132
rect 22465 41123 22523 41129
rect 22336 41092 22381 41120
rect 22336 41080 22342 41092
rect 22465 41089 22477 41123
rect 22511 41120 22523 41123
rect 23658 41120 23664 41132
rect 22511 41092 23664 41120
rect 22511 41089 22523 41092
rect 22465 41083 22523 41089
rect 23658 41080 23664 41092
rect 23716 41080 23722 41132
rect 24946 41120 24952 41132
rect 24907 41092 24952 41120
rect 24946 41080 24952 41092
rect 25004 41080 25010 41132
rect 25424 41129 25452 41160
rect 27706 41148 27712 41160
rect 27764 41148 27770 41200
rect 28644 41188 28672 41228
rect 28721 41225 28733 41259
rect 28767 41256 28779 41259
rect 29086 41256 29092 41268
rect 28767 41228 29092 41256
rect 28767 41225 28779 41228
rect 28721 41219 28779 41225
rect 29086 41216 29092 41228
rect 29144 41216 29150 41268
rect 29273 41259 29331 41265
rect 29273 41225 29285 41259
rect 29319 41256 29331 41259
rect 29914 41256 29920 41268
rect 29319 41228 29920 41256
rect 29319 41225 29331 41228
rect 29273 41219 29331 41225
rect 29914 41216 29920 41228
rect 29972 41216 29978 41268
rect 30650 41256 30656 41268
rect 30611 41228 30656 41256
rect 30650 41216 30656 41228
rect 30708 41216 30714 41268
rect 42334 41256 42340 41268
rect 31726 41228 42340 41256
rect 31726 41188 31754 41228
rect 42334 41216 42340 41228
rect 42392 41216 42398 41268
rect 42429 41259 42487 41265
rect 42429 41225 42441 41259
rect 42475 41256 42487 41259
rect 45738 41256 45744 41268
rect 42475 41228 45744 41256
rect 42475 41225 42487 41228
rect 42429 41219 42487 41225
rect 45738 41216 45744 41228
rect 45796 41216 45802 41268
rect 28644 41160 31754 41188
rect 35152 41191 35210 41197
rect 35152 41157 35164 41191
rect 35198 41188 35210 41191
rect 35250 41188 35256 41200
rect 35198 41160 35256 41188
rect 35198 41157 35210 41160
rect 35152 41151 35210 41157
rect 35250 41148 35256 41160
rect 35308 41148 35314 41200
rect 37550 41148 37556 41200
rect 37608 41188 37614 41200
rect 37608 41160 38148 41188
rect 37608 41148 37614 41160
rect 38120 41132 38148 41160
rect 39022 41148 39028 41200
rect 39080 41188 39086 41200
rect 39178 41191 39236 41197
rect 39178 41188 39190 41191
rect 39080 41160 39190 41188
rect 39080 41148 39086 41160
rect 39178 41157 39190 41160
rect 39224 41157 39236 41191
rect 39178 41151 39236 41157
rect 42518 41148 42524 41200
rect 42576 41188 42582 41200
rect 42886 41188 42892 41200
rect 42576 41160 42892 41188
rect 42576 41148 42582 41160
rect 42886 41148 42892 41160
rect 42944 41148 42950 41200
rect 45370 41148 45376 41200
rect 45428 41188 45434 41200
rect 45428 41160 46152 41188
rect 45428 41148 45434 41160
rect 25409 41123 25467 41129
rect 25409 41089 25421 41123
rect 25455 41089 25467 41123
rect 25409 41083 25467 41089
rect 27525 41123 27583 41129
rect 27525 41089 27537 41123
rect 27571 41089 27583 41123
rect 28442 41120 28448 41132
rect 28403 41092 28448 41120
rect 27525 41083 27583 41089
rect 21928 40956 22140 40984
rect 24394 40944 24400 40996
rect 24452 40984 24458 40996
rect 25501 40987 25559 40993
rect 25501 40984 25513 40987
rect 24452 40956 25513 40984
rect 24452 40944 24458 40956
rect 25501 40953 25513 40956
rect 25547 40953 25559 40987
rect 25501 40947 25559 40953
rect 27246 40944 27252 40996
rect 27304 40984 27310 40996
rect 27540 40984 27568 41083
rect 28442 41080 28448 41092
rect 28500 41080 28506 41132
rect 28537 41123 28595 41129
rect 28537 41089 28549 41123
rect 28583 41089 28595 41123
rect 28537 41083 28595 41089
rect 28258 41012 28264 41064
rect 28316 41052 28322 41064
rect 28552 41052 28580 41083
rect 29086 41080 29092 41132
rect 29144 41120 29150 41132
rect 29181 41123 29239 41129
rect 29181 41120 29193 41123
rect 29144 41092 29193 41120
rect 29144 41080 29150 41092
rect 29181 41089 29193 41092
rect 29227 41089 29239 41123
rect 30009 41123 30067 41129
rect 30009 41120 30021 41123
rect 29181 41083 29239 41089
rect 29288 41092 30021 41120
rect 29288 41052 29316 41092
rect 30009 41089 30021 41092
rect 30055 41089 30067 41123
rect 30009 41083 30067 41089
rect 30193 41123 30251 41129
rect 30193 41089 30205 41123
rect 30239 41120 30251 41123
rect 30837 41123 30895 41129
rect 30837 41120 30849 41123
rect 30239 41092 30849 41120
rect 30239 41089 30251 41092
rect 30193 41083 30251 41089
rect 30837 41089 30849 41092
rect 30883 41089 30895 41123
rect 32490 41120 32496 41132
rect 32451 41092 32496 41120
rect 30837 41083 30895 41089
rect 32490 41080 32496 41092
rect 32548 41080 32554 41132
rect 32674 41120 32680 41132
rect 32635 41092 32680 41120
rect 32674 41080 32680 41092
rect 32732 41080 32738 41132
rect 34422 41080 34428 41132
rect 34480 41120 34486 41132
rect 34885 41123 34943 41129
rect 34885 41120 34897 41123
rect 34480 41092 34897 41120
rect 34480 41080 34486 41092
rect 34885 41089 34897 41092
rect 34931 41089 34943 41123
rect 37274 41120 37280 41132
rect 37235 41092 37280 41120
rect 34885 41083 34943 41089
rect 37274 41080 37280 41092
rect 37332 41080 37338 41132
rect 37458 41120 37464 41132
rect 37419 41092 37464 41120
rect 37458 41080 37464 41092
rect 37516 41120 37522 41132
rect 37734 41120 37740 41132
rect 37516 41092 37740 41120
rect 37516 41080 37522 41092
rect 37734 41080 37740 41092
rect 37792 41080 37798 41132
rect 37826 41080 37832 41132
rect 37884 41080 37890 41132
rect 38102 41120 38108 41132
rect 38063 41092 38108 41120
rect 38102 41080 38108 41092
rect 38160 41080 38166 41132
rect 38378 41080 38384 41132
rect 38436 41120 38442 41132
rect 38933 41123 38991 41129
rect 38933 41120 38945 41123
rect 38436 41092 38945 41120
rect 38436 41080 38442 41092
rect 38933 41089 38945 41092
rect 38979 41089 38991 41123
rect 42705 41123 42763 41129
rect 42705 41120 42717 41123
rect 38933 41083 38991 41089
rect 40052 41092 42717 41120
rect 28316 41024 29316 41052
rect 29825 41055 29883 41061
rect 28316 41012 28322 41024
rect 29825 41021 29837 41055
rect 29871 41052 29883 41055
rect 31294 41052 31300 41064
rect 29871 41024 31300 41052
rect 29871 41021 29883 41024
rect 29825 41015 29883 41021
rect 31294 41012 31300 41024
rect 31352 41052 31358 41064
rect 33413 41055 33471 41061
rect 33413 41052 33425 41055
rect 31352 41024 33425 41052
rect 31352 41012 31358 41024
rect 33413 41021 33425 41024
rect 33459 41021 33471 41055
rect 33413 41015 33471 41021
rect 33502 41012 33508 41064
rect 33560 41061 33566 41064
rect 33560 41055 33588 41061
rect 33576 41021 33588 41055
rect 33560 41015 33588 41021
rect 33689 41055 33747 41061
rect 33689 41021 33701 41055
rect 33735 41052 33747 41055
rect 34514 41052 34520 41064
rect 33735 41024 34520 41052
rect 33735 41021 33747 41024
rect 33689 41015 33747 41021
rect 33560 41012 33566 41015
rect 34514 41012 34520 41024
rect 34572 41012 34578 41064
rect 37844 41052 37872 41080
rect 38654 41052 38660 41064
rect 37844 41024 38660 41052
rect 38654 41012 38660 41024
rect 38712 41012 38718 41064
rect 29086 40984 29092 40996
rect 27304 40956 29092 40984
rect 27304 40944 27310 40956
rect 29086 40944 29092 40956
rect 29144 40944 29150 40996
rect 33137 40987 33195 40993
rect 33137 40953 33149 40987
rect 33183 40953 33195 40987
rect 33137 40947 33195 40953
rect 24670 40876 24676 40928
rect 24728 40916 24734 40928
rect 24765 40919 24823 40925
rect 24765 40916 24777 40919
rect 24728 40888 24777 40916
rect 24728 40876 24734 40888
rect 24765 40885 24777 40888
rect 24811 40885 24823 40919
rect 24765 40879 24823 40885
rect 25866 40876 25872 40928
rect 25924 40916 25930 40928
rect 26050 40916 26056 40928
rect 25924 40888 26056 40916
rect 25924 40876 25930 40888
rect 26050 40876 26056 40888
rect 26108 40876 26114 40928
rect 28442 40876 28448 40928
rect 28500 40916 28506 40928
rect 28994 40916 29000 40928
rect 28500 40888 29000 40916
rect 28500 40876 28506 40888
rect 28994 40876 29000 40888
rect 29052 40876 29058 40928
rect 33152 40916 33180 40947
rect 37550 40944 37556 40996
rect 37608 40984 37614 40996
rect 38289 40987 38347 40993
rect 38289 40984 38301 40987
rect 37608 40956 38301 40984
rect 37608 40944 37614 40956
rect 38289 40953 38301 40956
rect 38335 40984 38347 40987
rect 38930 40984 38936 40996
rect 38335 40956 38936 40984
rect 38335 40953 38347 40956
rect 38289 40947 38347 40953
rect 38930 40944 38936 40956
rect 38988 40944 38994 40996
rect 33870 40916 33876 40928
rect 33152 40888 33876 40916
rect 33870 40876 33876 40888
rect 33928 40876 33934 40928
rect 34333 40919 34391 40925
rect 34333 40885 34345 40919
rect 34379 40916 34391 40919
rect 35526 40916 35532 40928
rect 34379 40888 35532 40916
rect 34379 40885 34391 40888
rect 34333 40879 34391 40885
rect 35526 40876 35532 40888
rect 35584 40876 35590 40928
rect 35618 40876 35624 40928
rect 35676 40916 35682 40928
rect 36265 40919 36323 40925
rect 36265 40916 36277 40919
rect 35676 40888 36277 40916
rect 35676 40876 35682 40888
rect 36265 40885 36277 40888
rect 36311 40885 36323 40919
rect 37642 40916 37648 40928
rect 37603 40888 37648 40916
rect 36265 40879 36323 40885
rect 37642 40876 37648 40888
rect 37700 40876 37706 40928
rect 38378 40876 38384 40928
rect 38436 40916 38442 40928
rect 40052 40916 40080 41092
rect 42705 41089 42717 41092
rect 42751 41089 42763 41123
rect 42705 41083 42763 41089
rect 43441 41123 43499 41129
rect 43441 41089 43453 41123
rect 43487 41089 43499 41123
rect 43441 41083 43499 41089
rect 40126 41012 40132 41064
rect 40184 41052 40190 41064
rect 41049 41055 41107 41061
rect 41049 41052 41061 41055
rect 40184 41024 41061 41052
rect 40184 41012 40190 41024
rect 41049 41021 41061 41024
rect 41095 41021 41107 41055
rect 41049 41015 41107 41021
rect 41325 41055 41383 41061
rect 41325 41021 41337 41055
rect 41371 41052 41383 41055
rect 41506 41052 41512 41064
rect 41371 41024 41512 41052
rect 41371 41021 41383 41024
rect 41325 41015 41383 41021
rect 41506 41012 41512 41024
rect 41564 41012 41570 41064
rect 42610 41052 42616 41064
rect 42571 41024 42616 41052
rect 42610 41012 42616 41024
rect 42668 41012 42674 41064
rect 42794 41052 42800 41064
rect 42755 41024 42800 41052
rect 42794 41012 42800 41024
rect 42852 41012 42858 41064
rect 42886 41012 42892 41064
rect 42944 41052 42950 41064
rect 43456 41052 43484 41083
rect 43898 41080 43904 41132
rect 43956 41120 43962 41132
rect 44361 41123 44419 41129
rect 44361 41120 44373 41123
rect 43956 41092 44373 41120
rect 43956 41080 43962 41092
rect 44361 41089 44373 41092
rect 44407 41089 44419 41123
rect 44361 41083 44419 41089
rect 45922 41080 45928 41132
rect 45980 41129 45986 41132
rect 46124 41129 46152 41160
rect 46290 41148 46296 41200
rect 46348 41148 46354 41200
rect 48866 41188 48872 41200
rect 48827 41160 48872 41188
rect 48866 41148 48872 41160
rect 48924 41148 48930 41200
rect 45980 41123 46029 41129
rect 45980 41089 45983 41123
rect 46017 41089 46029 41123
rect 45980 41083 46029 41089
rect 46109 41123 46167 41129
rect 46109 41089 46121 41123
rect 46155 41089 46167 41123
rect 46109 41083 46167 41089
rect 46201 41123 46259 41129
rect 46201 41089 46213 41123
rect 46247 41089 46259 41123
rect 46308 41120 46336 41148
rect 46385 41123 46443 41129
rect 46385 41120 46397 41123
rect 46308 41092 46397 41120
rect 46201 41083 46259 41089
rect 46385 41089 46397 41092
rect 46431 41089 46443 41123
rect 46385 41083 46443 41089
rect 45980 41080 45986 41083
rect 42944 41024 42989 41052
rect 43088 41024 43484 41052
rect 42944 41012 42950 41024
rect 40954 40944 40960 40996
rect 41012 40984 41018 40996
rect 43088 40984 43116 41024
rect 46216 40984 46244 41083
rect 67266 41080 67272 41132
rect 67324 41120 67330 41132
rect 67453 41123 67511 41129
rect 67453 41120 67465 41123
rect 67324 41092 67465 41120
rect 67324 41080 67330 41092
rect 67453 41089 67465 41092
rect 67499 41089 67511 41123
rect 67453 41083 67511 41089
rect 46290 41012 46296 41064
rect 46348 41052 46354 41064
rect 48038 41052 48044 41064
rect 46348 41024 48044 41052
rect 46348 41012 46354 41024
rect 48038 41012 48044 41024
rect 48096 41012 48102 41064
rect 48685 41055 48743 41061
rect 48685 41021 48697 41055
rect 48731 41021 48743 41055
rect 48685 41015 48743 41021
rect 50525 41055 50583 41061
rect 50525 41021 50537 41055
rect 50571 41052 50583 41055
rect 60734 41052 60740 41064
rect 50571 41024 60740 41052
rect 50571 41021 50583 41024
rect 50525 41015 50583 41021
rect 41012 40956 43116 40984
rect 43456 40956 46244 40984
rect 41012 40944 41018 40956
rect 40310 40916 40316 40928
rect 38436 40888 40080 40916
rect 40271 40888 40316 40916
rect 38436 40876 38442 40888
rect 40310 40876 40316 40888
rect 40368 40876 40374 40928
rect 41966 40876 41972 40928
rect 42024 40916 42030 40928
rect 43456 40916 43484 40956
rect 46382 40944 46388 40996
rect 46440 40984 46446 40996
rect 48700 40984 48728 41015
rect 60734 41012 60740 41024
rect 60792 41012 60798 41064
rect 46440 40956 48728 40984
rect 46440 40944 46446 40956
rect 43622 40916 43628 40928
rect 42024 40888 43484 40916
rect 43583 40888 43628 40916
rect 42024 40876 42030 40888
rect 43622 40876 43628 40888
rect 43680 40876 43686 40928
rect 44174 40916 44180 40928
rect 44135 40888 44180 40916
rect 44174 40876 44180 40888
rect 44232 40876 44238 40928
rect 45738 40916 45744 40928
rect 45699 40888 45744 40916
rect 45738 40876 45744 40888
rect 45796 40876 45802 40928
rect 66254 40876 66260 40928
rect 66312 40916 66318 40928
rect 66993 40919 67051 40925
rect 66993 40916 67005 40919
rect 66312 40888 67005 40916
rect 66312 40876 66318 40888
rect 66993 40885 67005 40888
rect 67039 40885 67051 40919
rect 66993 40879 67051 40885
rect 67082 40876 67088 40928
rect 67140 40916 67146 40928
rect 67545 40919 67603 40925
rect 67545 40916 67557 40919
rect 67140 40888 67557 40916
rect 67140 40876 67146 40888
rect 67545 40885 67557 40888
rect 67591 40885 67603 40919
rect 67545 40879 67603 40885
rect 1104 40826 68816 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 65654 40826
rect 65706 40774 65718 40826
rect 65770 40774 65782 40826
rect 65834 40774 65846 40826
rect 65898 40774 65910 40826
rect 65962 40774 68816 40826
rect 1104 40752 68816 40774
rect 22186 40712 22192 40724
rect 21928 40684 22192 40712
rect 6886 40616 19748 40644
rect 3234 40400 3240 40452
rect 3292 40440 3298 40452
rect 6886 40440 6914 40616
rect 19242 40576 19248 40588
rect 19203 40548 19248 40576
rect 19242 40536 19248 40548
rect 19300 40536 19306 40588
rect 19720 40585 19748 40616
rect 19705 40579 19763 40585
rect 19705 40545 19717 40579
rect 19751 40545 19763 40579
rect 19705 40539 19763 40545
rect 18509 40511 18567 40517
rect 18509 40477 18521 40511
rect 18555 40477 18567 40511
rect 18509 40471 18567 40477
rect 3292 40412 6914 40440
rect 3292 40400 3298 40412
rect 18524 40372 18552 40471
rect 21266 40468 21272 40520
rect 21324 40508 21330 40520
rect 21928 40517 21956 40684
rect 22186 40672 22192 40684
rect 22244 40712 22250 40724
rect 22738 40712 22744 40724
rect 22244 40684 22744 40712
rect 22244 40672 22250 40684
rect 22738 40672 22744 40684
rect 22796 40712 22802 40724
rect 22796 40684 31754 40712
rect 22796 40672 22802 40684
rect 22002 40604 22008 40656
rect 22060 40604 22066 40656
rect 27617 40647 27675 40653
rect 27617 40613 27629 40647
rect 27663 40613 27675 40647
rect 31726 40644 31754 40684
rect 34514 40672 34520 40724
rect 34572 40712 34578 40724
rect 34790 40712 34796 40724
rect 34572 40684 34796 40712
rect 34572 40672 34578 40684
rect 34790 40672 34796 40684
rect 34848 40672 34854 40724
rect 35342 40712 35348 40724
rect 35303 40684 35348 40712
rect 35342 40672 35348 40684
rect 35400 40672 35406 40724
rect 35434 40672 35440 40724
rect 35492 40712 35498 40724
rect 35529 40715 35587 40721
rect 35529 40712 35541 40715
rect 35492 40684 35541 40712
rect 35492 40672 35498 40684
rect 35529 40681 35541 40684
rect 35575 40681 35587 40715
rect 35529 40675 35587 40681
rect 36265 40715 36323 40721
rect 36265 40681 36277 40715
rect 36311 40712 36323 40715
rect 37826 40712 37832 40724
rect 36311 40684 37832 40712
rect 36311 40681 36323 40684
rect 36265 40675 36323 40681
rect 37826 40672 37832 40684
rect 37884 40672 37890 40724
rect 42610 40672 42616 40724
rect 42668 40712 42674 40724
rect 42889 40715 42947 40721
rect 42889 40712 42901 40715
rect 42668 40684 42901 40712
rect 42668 40672 42674 40684
rect 42889 40681 42901 40684
rect 42935 40681 42947 40715
rect 43898 40712 43904 40724
rect 43859 40684 43904 40712
rect 42889 40675 42947 40681
rect 43898 40672 43904 40684
rect 43956 40672 43962 40724
rect 48038 40712 48044 40724
rect 47999 40684 48044 40712
rect 48038 40672 48044 40684
rect 48096 40672 48102 40724
rect 37550 40644 37556 40656
rect 31726 40616 37556 40644
rect 27617 40607 27675 40613
rect 22020 40517 22048 40604
rect 23658 40576 23664 40588
rect 22204 40548 23664 40576
rect 22204 40517 22232 40548
rect 23658 40536 23664 40548
rect 23716 40536 23722 40588
rect 24394 40576 24400 40588
rect 24355 40548 24400 40576
rect 24394 40536 24400 40548
rect 24452 40536 24458 40588
rect 27632 40576 27660 40607
rect 37550 40604 37556 40616
rect 37608 40604 37614 40656
rect 37642 40604 37648 40656
rect 37700 40644 37706 40656
rect 41049 40647 41107 40653
rect 37700 40616 38608 40644
rect 37700 40604 37706 40616
rect 28074 40576 28080 40588
rect 27632 40548 28080 40576
rect 28074 40536 28080 40548
rect 28132 40536 28138 40588
rect 29270 40536 29276 40588
rect 29328 40576 29334 40588
rect 37274 40576 37280 40588
rect 29328 40548 37280 40576
rect 29328 40536 29334 40548
rect 37274 40536 37280 40548
rect 37332 40536 37338 40588
rect 38470 40576 38476 40588
rect 38431 40548 38476 40576
rect 38470 40536 38476 40548
rect 38528 40536 38534 40588
rect 38580 40585 38608 40616
rect 41049 40613 41061 40647
rect 41095 40644 41107 40647
rect 41414 40644 41420 40656
rect 41095 40616 41420 40644
rect 41095 40613 41107 40616
rect 41049 40607 41107 40613
rect 41414 40604 41420 40616
rect 41472 40604 41478 40656
rect 38565 40579 38623 40585
rect 38565 40545 38577 40579
rect 38611 40545 38623 40579
rect 38565 40539 38623 40545
rect 38657 40579 38715 40585
rect 38657 40545 38669 40579
rect 38703 40576 38715 40579
rect 39022 40576 39028 40588
rect 38703 40548 39028 40576
rect 38703 40545 38715 40548
rect 38657 40539 38715 40545
rect 39022 40536 39028 40548
rect 39080 40536 39086 40588
rect 42334 40536 42340 40588
rect 42392 40576 42398 40588
rect 45002 40576 45008 40588
rect 42392 40548 45008 40576
rect 42392 40536 42398 40548
rect 45002 40536 45008 40548
rect 45060 40576 45066 40588
rect 46658 40576 46664 40588
rect 45060 40548 45508 40576
rect 46619 40548 46664 40576
rect 45060 40536 45066 40548
rect 21775 40511 21833 40517
rect 21775 40508 21787 40511
rect 21324 40480 21787 40508
rect 21324 40468 21330 40480
rect 21775 40477 21787 40480
rect 21821 40477 21833 40511
rect 21775 40471 21833 40477
rect 21913 40511 21971 40517
rect 21913 40477 21925 40511
rect 21959 40477 21971 40511
rect 21913 40471 21971 40477
rect 22005 40511 22063 40517
rect 22005 40477 22017 40511
rect 22051 40477 22063 40511
rect 22005 40471 22063 40477
rect 22189 40511 22247 40517
rect 22189 40477 22201 40511
rect 22235 40477 22247 40511
rect 22189 40471 22247 40477
rect 23201 40511 23259 40517
rect 23201 40477 23213 40511
rect 23247 40508 23259 40511
rect 23290 40508 23296 40520
rect 23247 40480 23296 40508
rect 23247 40477 23259 40480
rect 23201 40471 23259 40477
rect 23290 40468 23296 40480
rect 23348 40468 23354 40520
rect 24670 40517 24676 40520
rect 24664 40508 24676 40517
rect 24631 40480 24676 40508
rect 24664 40471 24676 40480
rect 24670 40468 24676 40471
rect 24728 40468 24734 40520
rect 26234 40508 26240 40520
rect 26195 40480 26240 40508
rect 26234 40468 26240 40480
rect 26292 40468 26298 40520
rect 28258 40508 28264 40520
rect 28219 40480 28264 40508
rect 28258 40468 28264 40480
rect 28316 40468 28322 40520
rect 29086 40468 29092 40520
rect 29144 40508 29150 40520
rect 29549 40511 29607 40517
rect 29549 40508 29561 40511
rect 29144 40480 29561 40508
rect 29144 40468 29150 40480
rect 29549 40477 29561 40480
rect 29595 40477 29607 40511
rect 29549 40471 29607 40477
rect 33042 40468 33048 40520
rect 33100 40508 33106 40520
rect 36449 40511 36507 40517
rect 33100 40480 35756 40508
rect 33100 40468 33106 40480
rect 18601 40443 18659 40449
rect 18601 40409 18613 40443
rect 18647 40440 18659 40443
rect 19429 40443 19487 40449
rect 19429 40440 19441 40443
rect 18647 40412 19441 40440
rect 18647 40409 18659 40412
rect 18601 40403 18659 40409
rect 19429 40409 19441 40412
rect 19475 40409 19487 40443
rect 19429 40403 19487 40409
rect 26504 40443 26562 40449
rect 26504 40409 26516 40443
rect 26550 40440 26562 40443
rect 26970 40440 26976 40452
rect 26550 40412 26976 40440
rect 26550 40409 26562 40412
rect 26504 40403 26562 40409
rect 26970 40400 26976 40412
rect 27028 40400 27034 40452
rect 33502 40440 33508 40452
rect 27540 40412 33508 40440
rect 19978 40372 19984 40384
rect 18524 40344 19984 40372
rect 19978 40332 19984 40344
rect 20036 40332 20042 40384
rect 21542 40372 21548 40384
rect 21503 40344 21548 40372
rect 21542 40332 21548 40344
rect 21600 40332 21606 40384
rect 23382 40372 23388 40384
rect 23343 40344 23388 40372
rect 23382 40332 23388 40344
rect 23440 40332 23446 40384
rect 25130 40332 25136 40384
rect 25188 40372 25194 40384
rect 25777 40375 25835 40381
rect 25777 40372 25789 40375
rect 25188 40344 25789 40372
rect 25188 40332 25194 40344
rect 25777 40341 25789 40344
rect 25823 40372 25835 40375
rect 27540 40372 27568 40412
rect 33502 40400 33508 40412
rect 33560 40400 33566 40452
rect 35158 40440 35164 40452
rect 35071 40412 35164 40440
rect 35158 40400 35164 40412
rect 35216 40440 35222 40452
rect 35618 40440 35624 40452
rect 35216 40412 35624 40440
rect 35216 40400 35222 40412
rect 35618 40400 35624 40412
rect 35676 40400 35682 40452
rect 35728 40440 35756 40480
rect 36449 40477 36461 40511
rect 36495 40508 36507 40511
rect 37366 40508 37372 40520
rect 36495 40480 37372 40508
rect 36495 40477 36507 40480
rect 36449 40471 36507 40477
rect 37366 40468 37372 40480
rect 37424 40468 37430 40520
rect 38749 40511 38807 40517
rect 38749 40477 38761 40511
rect 38795 40508 38807 40511
rect 39114 40508 39120 40520
rect 38795 40480 39120 40508
rect 38795 40477 38807 40480
rect 38749 40471 38807 40477
rect 39114 40468 39120 40480
rect 39172 40508 39178 40520
rect 39390 40508 39396 40520
rect 39172 40480 39396 40508
rect 39172 40468 39178 40480
rect 39390 40468 39396 40480
rect 39448 40468 39454 40520
rect 41233 40511 41291 40517
rect 41233 40477 41245 40511
rect 41279 40477 41291 40511
rect 41233 40471 41291 40477
rect 43625 40511 43683 40517
rect 43625 40477 43637 40511
rect 43671 40477 43683 40511
rect 43625 40471 43683 40477
rect 37001 40443 37059 40449
rect 37001 40440 37013 40443
rect 35728 40412 37013 40440
rect 37001 40409 37013 40412
rect 37047 40440 37059 40443
rect 37734 40440 37740 40452
rect 37047 40412 37740 40440
rect 37047 40409 37059 40412
rect 37001 40403 37059 40409
rect 37734 40400 37740 40412
rect 37792 40400 37798 40452
rect 38654 40400 38660 40452
rect 38712 40440 38718 40452
rect 39758 40440 39764 40452
rect 38712 40412 39764 40440
rect 38712 40400 38718 40412
rect 39758 40400 39764 40412
rect 39816 40440 39822 40452
rect 41248 40440 41276 40471
rect 42518 40440 42524 40452
rect 39816 40412 41276 40440
rect 42479 40412 42524 40440
rect 39816 40400 39822 40412
rect 42518 40400 42524 40412
rect 42576 40400 42582 40452
rect 42705 40443 42763 40449
rect 42705 40409 42717 40443
rect 42751 40440 42763 40443
rect 43640 40440 43668 40471
rect 43714 40468 43720 40520
rect 43772 40508 43778 40520
rect 45480 40517 45508 40548
rect 46658 40536 46664 40548
rect 46716 40536 46722 40588
rect 66254 40576 66260 40588
rect 66215 40548 66260 40576
rect 66254 40536 66260 40548
rect 66312 40536 66318 40588
rect 66441 40579 66499 40585
rect 66441 40545 66453 40579
rect 66487 40576 66499 40579
rect 67082 40576 67088 40588
rect 66487 40548 67088 40576
rect 66487 40545 66499 40548
rect 66441 40539 66499 40545
rect 67082 40536 67088 40548
rect 67140 40536 67146 40588
rect 68094 40576 68100 40588
rect 68055 40548 68100 40576
rect 68094 40536 68100 40548
rect 68152 40536 68158 40588
rect 45465 40511 45523 40517
rect 43772 40480 43817 40508
rect 43772 40468 43778 40480
rect 45465 40477 45477 40511
rect 45511 40477 45523 40511
rect 45465 40471 45523 40477
rect 45738 40468 45744 40520
rect 45796 40508 45802 40520
rect 46917 40511 46975 40517
rect 46917 40508 46929 40511
rect 45796 40480 46929 40508
rect 45796 40468 45802 40480
rect 46917 40477 46929 40480
rect 46963 40477 46975 40511
rect 48774 40508 48780 40520
rect 48735 40480 48780 40508
rect 46917 40471 46975 40477
rect 48774 40468 48780 40480
rect 48832 40468 48838 40520
rect 45186 40440 45192 40452
rect 42751 40412 45192 40440
rect 42751 40409 42763 40412
rect 42705 40403 42763 40409
rect 45186 40400 45192 40412
rect 45244 40400 45250 40452
rect 28442 40372 28448 40384
rect 25823 40344 27568 40372
rect 28403 40344 28448 40372
rect 25823 40341 25835 40344
rect 25777 40335 25835 40341
rect 28442 40332 28448 40344
rect 28500 40332 28506 40384
rect 29270 40332 29276 40384
rect 29328 40372 29334 40384
rect 29733 40375 29791 40381
rect 29733 40372 29745 40375
rect 29328 40344 29745 40372
rect 29328 40332 29334 40344
rect 29733 40341 29745 40344
rect 29779 40341 29791 40375
rect 29733 40335 29791 40341
rect 34698 40332 34704 40384
rect 34756 40372 34762 40384
rect 35342 40372 35348 40384
rect 35400 40381 35406 40384
rect 35400 40375 35419 40381
rect 34756 40344 35348 40372
rect 34756 40332 34762 40344
rect 35342 40332 35348 40344
rect 35407 40341 35419 40375
rect 35400 40335 35419 40341
rect 37277 40375 37335 40381
rect 37277 40341 37289 40375
rect 37323 40372 37335 40375
rect 38010 40372 38016 40384
rect 37323 40344 38016 40372
rect 37323 40341 37335 40344
rect 37277 40335 37335 40341
rect 35400 40332 35406 40335
rect 38010 40332 38016 40344
rect 38068 40332 38074 40384
rect 38289 40375 38347 40381
rect 38289 40341 38301 40375
rect 38335 40372 38347 40375
rect 38746 40372 38752 40384
rect 38335 40344 38752 40372
rect 38335 40341 38347 40344
rect 38289 40335 38347 40341
rect 38746 40332 38752 40344
rect 38804 40332 38810 40384
rect 45649 40375 45707 40381
rect 45649 40341 45661 40375
rect 45695 40372 45707 40375
rect 46106 40372 46112 40384
rect 45695 40344 46112 40372
rect 45695 40341 45707 40344
rect 45649 40335 45707 40341
rect 46106 40332 46112 40344
rect 46164 40332 46170 40384
rect 48869 40375 48927 40381
rect 48869 40341 48881 40375
rect 48915 40372 48927 40375
rect 48958 40372 48964 40384
rect 48915 40344 48964 40372
rect 48915 40341 48927 40344
rect 48869 40335 48927 40341
rect 48958 40332 48964 40344
rect 49016 40332 49022 40384
rect 1104 40282 68816 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 68816 40282
rect 1104 40208 68816 40230
rect 22462 40168 22468 40180
rect 19936 40140 22468 40168
rect 19936 40100 19964 40140
rect 22462 40128 22468 40140
rect 22520 40128 22526 40180
rect 24946 40128 24952 40180
rect 25004 40168 25010 40180
rect 25409 40171 25467 40177
rect 25409 40168 25421 40171
rect 25004 40140 25421 40168
rect 25004 40128 25010 40140
rect 25409 40137 25421 40140
rect 25455 40137 25467 40171
rect 25409 40131 25467 40137
rect 26234 40128 26240 40180
rect 26292 40168 26298 40180
rect 26329 40171 26387 40177
rect 26329 40168 26341 40171
rect 26292 40140 26341 40168
rect 26292 40128 26298 40140
rect 26329 40137 26341 40140
rect 26375 40137 26387 40171
rect 26970 40168 26976 40180
rect 26931 40140 26976 40168
rect 26329 40131 26387 40137
rect 26970 40128 26976 40140
rect 27028 40128 27034 40180
rect 35158 40168 35164 40180
rect 33428 40140 35164 40168
rect 23382 40100 23388 40112
rect 19904 40072 19964 40100
rect 19996 40072 23388 40100
rect 19904 40041 19932 40072
rect 19996 40044 20024 40072
rect 19889 40035 19947 40041
rect 19889 40001 19901 40035
rect 19935 40001 19947 40035
rect 19889 39995 19947 40001
rect 19978 39992 19984 40044
rect 20036 39992 20042 40044
rect 20156 40035 20214 40041
rect 20156 40001 20168 40035
rect 20202 40032 20214 40035
rect 21542 40032 21548 40044
rect 20202 40004 21548 40032
rect 20202 40001 20214 40004
rect 20156 39995 20214 40001
rect 21542 39992 21548 40004
rect 21600 39992 21606 40044
rect 22664 40041 22692 40072
rect 23382 40060 23388 40072
rect 23440 40060 23446 40112
rect 28442 40100 28448 40112
rect 27172 40072 28448 40100
rect 22649 40035 22707 40041
rect 22649 40001 22661 40035
rect 22695 40001 22707 40035
rect 22649 39995 22707 40001
rect 22741 40035 22799 40041
rect 22741 40001 22753 40035
rect 22787 40032 22799 40035
rect 22830 40032 22836 40044
rect 22787 40004 22836 40032
rect 22787 40001 22799 40004
rect 22741 39995 22799 40001
rect 22830 39992 22836 40004
rect 22888 39992 22894 40044
rect 25130 40032 25136 40044
rect 25091 40004 25136 40032
rect 25130 39992 25136 40004
rect 25188 39992 25194 40044
rect 25222 39992 25228 40044
rect 25280 40032 25286 40044
rect 26326 40032 26332 40044
rect 25280 40004 25325 40032
rect 26287 40004 26332 40032
rect 25280 39992 25286 40004
rect 26326 39992 26332 40004
rect 26384 39992 26390 40044
rect 27172 40041 27200 40072
rect 28442 40060 28448 40072
rect 28500 40060 28506 40112
rect 32493 40103 32551 40109
rect 32493 40100 32505 40103
rect 31588 40072 32505 40100
rect 27157 40035 27215 40041
rect 27157 40001 27169 40035
rect 27203 40001 27215 40035
rect 28258 40032 28264 40044
rect 28219 40004 28264 40032
rect 27157 39995 27215 40001
rect 28258 39992 28264 40004
rect 28316 39992 28322 40044
rect 29270 40032 29276 40044
rect 29231 40004 29276 40032
rect 29270 39992 29276 40004
rect 29328 39992 29334 40044
rect 29540 40035 29598 40041
rect 29540 40001 29552 40035
rect 29586 40032 29598 40035
rect 30466 40032 30472 40044
rect 29586 40004 30472 40032
rect 29586 40001 29598 40004
rect 29540 39995 29598 40001
rect 30466 39992 30472 40004
rect 30524 39992 30530 40044
rect 31588 40041 31616 40072
rect 32493 40069 32505 40072
rect 32539 40069 32551 40103
rect 32493 40063 32551 40069
rect 31573 40035 31631 40041
rect 31573 40001 31585 40035
rect 31619 40001 31631 40035
rect 32306 40032 32312 40044
rect 32267 40004 32312 40032
rect 31573 39995 31631 40001
rect 32306 39992 32312 40004
rect 32364 39992 32370 40044
rect 33226 40032 33232 40044
rect 33187 40004 33232 40032
rect 33226 39992 33232 40004
rect 33284 39992 33290 40044
rect 33428 40041 33456 40140
rect 35158 40128 35164 40140
rect 35216 40128 35222 40180
rect 38102 40128 38108 40180
rect 38160 40168 38166 40180
rect 44358 40168 44364 40180
rect 38160 40140 44364 40168
rect 38160 40128 38166 40140
rect 44358 40128 44364 40140
rect 44416 40128 44422 40180
rect 45186 40168 45192 40180
rect 45147 40140 45192 40168
rect 45186 40128 45192 40140
rect 45244 40128 45250 40180
rect 46290 40128 46296 40180
rect 46348 40168 46354 40180
rect 46348 40140 46934 40168
rect 46348 40128 46354 40140
rect 37277 40103 37335 40109
rect 37277 40100 37289 40103
rect 36188 40072 37289 40100
rect 33413 40035 33471 40041
rect 33413 40001 33425 40035
rect 33459 40001 33471 40035
rect 33413 39995 33471 40001
rect 35069 40035 35127 40041
rect 35069 40001 35081 40035
rect 35115 40032 35127 40035
rect 36188 40032 36216 40072
rect 37277 40069 37289 40072
rect 37323 40069 37335 40103
rect 38194 40100 38200 40112
rect 38155 40072 38200 40100
rect 37277 40063 37335 40069
rect 38194 40060 38200 40072
rect 38252 40060 38258 40112
rect 39025 40103 39083 40109
rect 39025 40069 39037 40103
rect 39071 40100 39083 40103
rect 39206 40100 39212 40112
rect 39071 40072 39212 40100
rect 39071 40069 39083 40072
rect 39025 40063 39083 40069
rect 39206 40060 39212 40072
rect 39264 40100 39270 40112
rect 39574 40100 39580 40112
rect 39264 40072 39580 40100
rect 39264 40060 39270 40072
rect 39574 40060 39580 40072
rect 39632 40060 39638 40112
rect 41414 40060 41420 40112
rect 41472 40100 41478 40112
rect 42518 40100 42524 40112
rect 41472 40072 42524 40100
rect 41472 40060 41478 40072
rect 42518 40060 42524 40072
rect 42576 40060 42582 40112
rect 42705 40103 42763 40109
rect 42705 40069 42717 40103
rect 42751 40100 42763 40103
rect 43346 40100 43352 40112
rect 42751 40072 43352 40100
rect 42751 40069 42763 40072
rect 42705 40063 42763 40069
rect 43346 40060 43352 40072
rect 43404 40060 43410 40112
rect 44174 40060 44180 40112
rect 44232 40060 44238 40112
rect 46906 40100 46934 40140
rect 48130 40100 48136 40112
rect 46906 40072 48136 40100
rect 48130 40060 48136 40072
rect 48188 40060 48194 40112
rect 48958 40100 48964 40112
rect 48919 40072 48964 40100
rect 48958 40060 48964 40072
rect 49016 40060 49022 40112
rect 50617 40103 50675 40109
rect 50617 40069 50629 40103
rect 50663 40100 50675 40103
rect 66070 40100 66076 40112
rect 50663 40072 66076 40100
rect 50663 40069 50675 40072
rect 50617 40063 50675 40069
rect 66070 40060 66076 40072
rect 66128 40060 66134 40112
rect 67266 40100 67272 40112
rect 67227 40072 67272 40100
rect 67266 40060 67272 40072
rect 67324 40060 67330 40112
rect 35115 40004 36216 40032
rect 37461 40035 37519 40041
rect 35115 40001 35127 40004
rect 35069 39995 35127 40001
rect 37461 40001 37473 40035
rect 37507 40032 37519 40035
rect 37826 40032 37832 40044
rect 37507 40004 37832 40032
rect 37507 40001 37519 40004
rect 37461 39995 37519 40001
rect 37826 39992 37832 40004
rect 37884 39992 37890 40044
rect 40212 40035 40270 40041
rect 40212 40001 40224 40035
rect 40258 40032 40270 40035
rect 40494 40032 40500 40044
rect 40258 40004 40500 40032
rect 40258 40001 40270 40004
rect 40212 39995 40270 40001
rect 40494 39992 40500 40004
rect 40552 39992 40558 40044
rect 43622 39992 43628 40044
rect 43680 40032 43686 40044
rect 43809 40035 43867 40041
rect 43809 40032 43821 40035
rect 43680 40004 43821 40032
rect 43680 39992 43686 40004
rect 43809 40001 43821 40004
rect 43855 40001 43867 40035
rect 43809 39995 43867 40001
rect 44076 40035 44134 40041
rect 44076 40001 44088 40035
rect 44122 40032 44134 40035
rect 44192 40032 44220 40060
rect 44122 40004 44220 40032
rect 44122 40001 44134 40004
rect 44076 39995 44134 40001
rect 46290 39992 46296 40044
rect 46348 40041 46354 40044
rect 46348 40035 46397 40041
rect 46348 40001 46351 40035
rect 46385 40001 46397 40035
rect 46348 39995 46397 40001
rect 46477 40035 46535 40041
rect 46477 40001 46489 40035
rect 46523 40001 46535 40035
rect 46477 39995 46535 40001
rect 46348 39992 46354 39995
rect 27798 39924 27804 39976
rect 27856 39964 27862 39976
rect 27985 39967 28043 39973
rect 27985 39964 27997 39967
rect 27856 39936 27997 39964
rect 27856 39924 27862 39936
rect 27985 39933 27997 39936
rect 28031 39933 28043 39967
rect 27985 39927 28043 39933
rect 32125 39967 32183 39973
rect 32125 39933 32137 39967
rect 32171 39964 32183 39967
rect 32674 39964 32680 39976
rect 32171 39936 32680 39964
rect 32171 39933 32183 39936
rect 32125 39927 32183 39933
rect 32674 39924 32680 39936
rect 32732 39924 32738 39976
rect 34149 39967 34207 39973
rect 34149 39964 34161 39967
rect 32968 39936 34161 39964
rect 32968 39896 32996 39936
rect 34149 39933 34161 39936
rect 34195 39933 34207 39967
rect 34149 39927 34207 39933
rect 34238 39924 34244 39976
rect 34296 39973 34302 39976
rect 34296 39967 34324 39973
rect 34312 39933 34324 39967
rect 34296 39927 34324 39933
rect 34425 39967 34483 39973
rect 34425 39933 34437 39967
rect 34471 39964 34483 39967
rect 34790 39964 34796 39976
rect 34471 39936 34796 39964
rect 34471 39933 34483 39936
rect 34425 39927 34483 39933
rect 34296 39924 34302 39927
rect 34790 39924 34796 39936
rect 34848 39924 34854 39976
rect 39942 39964 39948 39976
rect 39903 39936 39948 39964
rect 39942 39924 39948 39936
rect 40000 39924 40006 39976
rect 30668 39868 32996 39896
rect 1394 39788 1400 39840
rect 1452 39828 1458 39840
rect 1673 39831 1731 39837
rect 1673 39828 1685 39831
rect 1452 39800 1685 39828
rect 1452 39788 1458 39800
rect 1673 39797 1685 39800
rect 1719 39797 1731 39831
rect 21266 39828 21272 39840
rect 21227 39800 21272 39828
rect 1673 39791 1731 39797
rect 21266 39788 21272 39800
rect 21324 39788 21330 39840
rect 30558 39788 30564 39840
rect 30616 39828 30622 39840
rect 30668 39837 30696 39868
rect 33226 39856 33232 39908
rect 33284 39896 33290 39908
rect 33594 39896 33600 39908
rect 33284 39868 33600 39896
rect 33284 39856 33290 39868
rect 33594 39856 33600 39868
rect 33652 39856 33658 39908
rect 33870 39896 33876 39908
rect 33831 39868 33876 39896
rect 33870 39856 33876 39868
rect 33928 39856 33934 39908
rect 37918 39856 37924 39908
rect 37976 39896 37982 39908
rect 38378 39896 38384 39908
rect 37976 39868 38384 39896
rect 37976 39856 37982 39868
rect 38378 39856 38384 39868
rect 38436 39856 38442 39908
rect 45370 39856 45376 39908
rect 45428 39896 45434 39908
rect 46492 39896 46520 39995
rect 46566 39992 46572 40044
rect 46624 40032 46630 40044
rect 46624 40004 46666 40032
rect 46624 39992 46630 40004
rect 46750 39992 46756 40044
rect 46808 40032 46814 40044
rect 48148 40032 48176 40060
rect 48777 40035 48835 40041
rect 48777 40032 48789 40035
rect 46808 40004 46853 40032
rect 48148 40004 48789 40032
rect 46808 39992 46814 40004
rect 48777 40001 48789 40004
rect 48823 40001 48835 40035
rect 48777 39995 48835 40001
rect 45428 39868 46520 39896
rect 45428 39856 45434 39868
rect 30653 39831 30711 39837
rect 30653 39828 30665 39831
rect 30616 39800 30665 39828
rect 30616 39788 30622 39800
rect 30653 39797 30665 39800
rect 30699 39797 30711 39831
rect 31386 39828 31392 39840
rect 31347 39800 31392 39828
rect 30653 39791 30711 39797
rect 31386 39788 31392 39800
rect 31444 39788 31450 39840
rect 37642 39828 37648 39840
rect 37603 39800 37648 39828
rect 37642 39788 37648 39800
rect 37700 39788 37706 39840
rect 39114 39828 39120 39840
rect 39075 39800 39120 39828
rect 39114 39788 39120 39800
rect 39172 39788 39178 39840
rect 41046 39788 41052 39840
rect 41104 39828 41110 39840
rect 41325 39831 41383 39837
rect 41325 39828 41337 39831
rect 41104 39800 41337 39828
rect 41104 39788 41110 39800
rect 41325 39797 41337 39800
rect 41371 39797 41383 39831
rect 41325 39791 41383 39797
rect 42610 39788 42616 39840
rect 42668 39828 42674 39840
rect 42889 39831 42947 39837
rect 42889 39828 42901 39831
rect 42668 39800 42901 39828
rect 42668 39788 42674 39800
rect 42889 39797 42901 39800
rect 42935 39797 42947 39831
rect 42889 39791 42947 39797
rect 46109 39831 46167 39837
rect 46109 39797 46121 39831
rect 46155 39828 46167 39831
rect 46842 39828 46848 39840
rect 46155 39800 46848 39828
rect 46155 39797 46167 39800
rect 46109 39791 46167 39797
rect 46842 39788 46848 39800
rect 46900 39788 46906 39840
rect 67358 39828 67364 39840
rect 67319 39800 67364 39828
rect 67358 39788 67364 39800
rect 67416 39788 67422 39840
rect 1104 39738 68816 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 65654 39738
rect 65706 39686 65718 39738
rect 65770 39686 65782 39738
rect 65834 39686 65846 39738
rect 65898 39686 65910 39738
rect 65962 39686 68816 39738
rect 1104 39664 68816 39686
rect 25774 39624 25780 39636
rect 25687 39596 25780 39624
rect 25774 39584 25780 39596
rect 25832 39624 25838 39636
rect 26142 39624 26148 39636
rect 25832 39596 26148 39624
rect 25832 39584 25838 39596
rect 26142 39584 26148 39596
rect 26200 39584 26206 39636
rect 26326 39584 26332 39636
rect 26384 39624 26390 39636
rect 26513 39627 26571 39633
rect 26513 39624 26525 39627
rect 26384 39596 26525 39624
rect 26384 39584 26390 39596
rect 26513 39593 26525 39596
rect 26559 39624 26571 39627
rect 27246 39624 27252 39636
rect 26559 39596 27252 39624
rect 26559 39593 26571 39596
rect 26513 39587 26571 39593
rect 27246 39584 27252 39596
rect 27304 39584 27310 39636
rect 30466 39624 30472 39636
rect 30427 39596 30472 39624
rect 30466 39584 30472 39596
rect 30524 39584 30530 39636
rect 32674 39624 32680 39636
rect 32587 39596 32680 39624
rect 32674 39584 32680 39596
rect 32732 39624 32738 39636
rect 34238 39624 34244 39636
rect 32732 39596 34244 39624
rect 32732 39584 32738 39596
rect 34238 39584 34244 39596
rect 34296 39584 34302 39636
rect 35345 39627 35403 39633
rect 35345 39593 35357 39627
rect 35391 39624 35403 39627
rect 35434 39624 35440 39636
rect 35391 39596 35440 39624
rect 35391 39593 35403 39596
rect 35345 39587 35403 39593
rect 35434 39584 35440 39596
rect 35492 39584 35498 39636
rect 39942 39584 39948 39636
rect 40000 39624 40006 39636
rect 40221 39627 40279 39633
rect 40221 39624 40233 39627
rect 40000 39596 40233 39624
rect 40000 39584 40006 39596
rect 40221 39593 40233 39596
rect 40267 39593 40279 39627
rect 40221 39587 40279 39593
rect 42429 39627 42487 39633
rect 42429 39593 42441 39627
rect 42475 39624 42487 39627
rect 46566 39624 46572 39636
rect 42475 39596 46572 39624
rect 42475 39593 42487 39596
rect 42429 39587 42487 39593
rect 46566 39584 46572 39596
rect 46624 39584 46630 39636
rect 48130 39624 48136 39636
rect 48091 39596 48136 39624
rect 48130 39584 48136 39596
rect 48188 39584 48194 39636
rect 29822 39556 29828 39568
rect 26804 39528 29828 39556
rect 1394 39488 1400 39500
rect 1355 39460 1400 39488
rect 1394 39448 1400 39460
rect 1452 39448 1458 39500
rect 2774 39488 2780 39500
rect 2735 39460 2780 39488
rect 2774 39448 2780 39460
rect 2832 39448 2838 39500
rect 19337 39491 19395 39497
rect 19337 39457 19349 39491
rect 19383 39488 19395 39491
rect 21266 39488 21272 39500
rect 19383 39460 21272 39488
rect 19383 39457 19395 39460
rect 19337 39451 19395 39457
rect 21266 39448 21272 39460
rect 21324 39448 21330 39500
rect 22462 39488 22468 39500
rect 22423 39460 22468 39488
rect 22462 39448 22468 39460
rect 22520 39448 22526 39500
rect 26804 39432 26832 39528
rect 29822 39516 29828 39528
rect 29880 39516 29886 39568
rect 37642 39516 37648 39568
rect 37700 39556 37706 39568
rect 37700 39528 41414 39556
rect 37700 39516 37706 39528
rect 29641 39491 29699 39497
rect 29641 39457 29653 39491
rect 29687 39488 29699 39491
rect 30558 39488 30564 39500
rect 29687 39460 30564 39488
rect 29687 39457 29699 39460
rect 29641 39451 29699 39457
rect 30558 39448 30564 39460
rect 30616 39448 30622 39500
rect 38838 39488 38844 39500
rect 38672 39460 38844 39488
rect 26329 39423 26387 39429
rect 26329 39389 26341 39423
rect 26375 39420 26387 39423
rect 26786 39420 26792 39432
rect 26375 39392 26792 39420
rect 26375 39389 26387 39392
rect 26329 39383 26387 39389
rect 26786 39380 26792 39392
rect 26844 39380 26850 39432
rect 27246 39420 27252 39432
rect 27207 39392 27252 39420
rect 27246 39380 27252 39392
rect 27304 39380 27310 39432
rect 28166 39420 28172 39432
rect 28127 39392 28172 39420
rect 28166 39380 28172 39392
rect 28224 39380 28230 39432
rect 28258 39380 28264 39432
rect 28316 39420 28322 39432
rect 29825 39423 29883 39429
rect 29825 39420 29837 39423
rect 28316 39392 29837 39420
rect 28316 39380 28322 39392
rect 29825 39389 29837 39392
rect 29871 39389 29883 39423
rect 29825 39383 29883 39389
rect 30009 39423 30067 39429
rect 30009 39389 30021 39423
rect 30055 39420 30067 39423
rect 30653 39423 30711 39429
rect 30653 39420 30665 39423
rect 30055 39392 30665 39420
rect 30055 39389 30067 39392
rect 30009 39383 30067 39389
rect 30653 39389 30665 39392
rect 30699 39389 30711 39423
rect 30653 39383 30711 39389
rect 31018 39380 31024 39432
rect 31076 39420 31082 39432
rect 31297 39423 31355 39429
rect 31297 39420 31309 39423
rect 31076 39392 31309 39420
rect 31076 39380 31082 39392
rect 31297 39389 31309 39392
rect 31343 39389 31355 39423
rect 31297 39383 31355 39389
rect 31386 39380 31392 39432
rect 31444 39420 31450 39432
rect 31553 39423 31611 39429
rect 31553 39420 31565 39423
rect 31444 39392 31565 39420
rect 31444 39380 31450 39392
rect 31553 39389 31565 39392
rect 31599 39389 31611 39423
rect 35434 39420 35440 39432
rect 31553 39383 31611 39389
rect 35176 39392 35440 39420
rect 1581 39355 1639 39361
rect 1581 39321 1593 39355
rect 1627 39352 1639 39355
rect 1854 39352 1860 39364
rect 1627 39324 1860 39352
rect 1627 39321 1639 39324
rect 1581 39315 1639 39321
rect 1854 39312 1860 39324
rect 1912 39312 1918 39364
rect 19521 39355 19579 39361
rect 19521 39321 19533 39355
rect 19567 39321 19579 39355
rect 19521 39315 19579 39321
rect 19426 39244 19432 39296
rect 19484 39284 19490 39296
rect 19536 39284 19564 39315
rect 20714 39312 20720 39364
rect 20772 39352 20778 39364
rect 21177 39355 21235 39361
rect 21177 39352 21189 39355
rect 20772 39324 21189 39352
rect 20772 39312 20778 39324
rect 21177 39321 21189 39324
rect 21223 39321 21235 39355
rect 21177 39315 21235 39321
rect 22554 39312 22560 39364
rect 22612 39352 22618 39364
rect 22710 39355 22768 39361
rect 22710 39352 22722 39355
rect 22612 39324 22722 39352
rect 22612 39312 22618 39324
rect 22710 39321 22722 39324
rect 22756 39321 22768 39355
rect 22710 39315 22768 39321
rect 25501 39355 25559 39361
rect 25501 39321 25513 39355
rect 25547 39352 25559 39355
rect 25866 39352 25872 39364
rect 25547 39324 25872 39352
rect 25547 39321 25559 39324
rect 25501 39315 25559 39321
rect 25866 39312 25872 39324
rect 25924 39312 25930 39364
rect 33594 39312 33600 39364
rect 33652 39352 33658 39364
rect 35176 39361 35204 39392
rect 35434 39380 35440 39392
rect 35492 39380 35498 39432
rect 37461 39423 37519 39429
rect 37461 39389 37473 39423
rect 37507 39420 37519 39423
rect 37826 39420 37832 39432
rect 37507 39392 37832 39420
rect 37507 39389 37519 39392
rect 37461 39383 37519 39389
rect 37826 39380 37832 39392
rect 37884 39380 37890 39432
rect 38470 39380 38476 39432
rect 38528 39416 38534 39432
rect 38672 39429 38700 39460
rect 38838 39448 38844 39460
rect 38896 39488 38902 39500
rect 40034 39488 40040 39500
rect 38896 39460 40040 39488
rect 38896 39448 38902 39460
rect 40034 39448 40040 39460
rect 40092 39448 40098 39500
rect 41386 39488 41414 39528
rect 45370 39516 45376 39568
rect 45428 39516 45434 39568
rect 42705 39491 42763 39497
rect 42705 39488 42717 39491
rect 41386 39460 42717 39488
rect 42705 39457 42717 39460
rect 42751 39457 42763 39491
rect 42886 39488 42892 39500
rect 42847 39460 42892 39488
rect 42705 39451 42763 39457
rect 42886 39448 42892 39460
rect 42944 39448 42950 39500
rect 38565 39423 38623 39429
rect 38565 39416 38577 39423
rect 38528 39389 38577 39416
rect 38611 39389 38623 39423
rect 38528 39388 38623 39389
rect 38528 39380 38534 39388
rect 38565 39383 38623 39388
rect 38654 39423 38712 39429
rect 38654 39389 38666 39423
rect 38700 39389 38712 39423
rect 38654 39383 38712 39389
rect 38746 39380 38752 39432
rect 38804 39420 38810 39432
rect 38933 39423 38991 39429
rect 38804 39392 38849 39420
rect 38804 39380 38810 39392
rect 38933 39389 38945 39423
rect 38979 39420 38991 39423
rect 39482 39420 39488 39432
rect 38979 39392 39488 39420
rect 38979 39389 38991 39392
rect 38933 39383 38991 39389
rect 39482 39380 39488 39392
rect 39540 39420 39546 39432
rect 39850 39420 39856 39432
rect 39540 39392 39856 39420
rect 39540 39380 39546 39392
rect 39850 39380 39856 39392
rect 39908 39380 39914 39432
rect 40405 39423 40463 39429
rect 40405 39389 40417 39423
rect 40451 39420 40463 39423
rect 40862 39420 40868 39432
rect 40451 39392 40868 39420
rect 40451 39389 40463 39392
rect 40405 39383 40463 39389
rect 40862 39380 40868 39392
rect 40920 39380 40926 39432
rect 41046 39420 41052 39432
rect 41007 39392 41052 39420
rect 41046 39380 41052 39392
rect 41104 39380 41110 39432
rect 41141 39423 41199 39429
rect 41141 39389 41153 39423
rect 41187 39420 41199 39423
rect 42610 39420 42616 39432
rect 41187 39392 42472 39420
rect 42571 39392 42616 39420
rect 41187 39389 41199 39392
rect 41141 39383 41199 39389
rect 35161 39355 35219 39361
rect 35161 39352 35173 39355
rect 33652 39324 35173 39352
rect 33652 39312 33658 39324
rect 35161 39321 35173 39324
rect 35207 39321 35219 39355
rect 35161 39315 35219 39321
rect 35250 39312 35256 39364
rect 35308 39352 35314 39364
rect 37277 39355 37335 39361
rect 37277 39352 37289 39355
rect 35308 39324 37289 39352
rect 35308 39312 35314 39324
rect 37277 39321 37289 39324
rect 37323 39321 37335 39355
rect 37277 39315 37335 39321
rect 37645 39355 37703 39361
rect 37645 39321 37657 39355
rect 37691 39352 37703 39355
rect 42334 39352 42340 39364
rect 37691 39324 38608 39352
rect 37691 39321 37703 39324
rect 37645 39315 37703 39321
rect 19484 39256 19564 39284
rect 19484 39244 19490 39256
rect 23750 39244 23756 39296
rect 23808 39284 23814 39296
rect 23845 39287 23903 39293
rect 23845 39284 23857 39287
rect 23808 39256 23857 39284
rect 23808 39244 23814 39256
rect 23845 39253 23857 39256
rect 23891 39253 23903 39287
rect 23845 39247 23903 39253
rect 27062 39244 27068 39296
rect 27120 39284 27126 39296
rect 27249 39287 27307 39293
rect 27249 39284 27261 39287
rect 27120 39256 27261 39284
rect 27120 39244 27126 39256
rect 27249 39253 27261 39256
rect 27295 39253 27307 39287
rect 27249 39247 27307 39253
rect 27890 39244 27896 39296
rect 27948 39284 27954 39296
rect 28445 39287 28503 39293
rect 28445 39284 28457 39287
rect 27948 39256 28457 39284
rect 27948 39244 27954 39256
rect 28445 39253 28457 39256
rect 28491 39253 28503 39287
rect 28445 39247 28503 39253
rect 35342 39244 35348 39296
rect 35400 39293 35406 39296
rect 35400 39287 35419 39293
rect 35407 39253 35419 39287
rect 35400 39247 35419 39253
rect 35529 39287 35587 39293
rect 35529 39253 35541 39287
rect 35575 39284 35587 39287
rect 36722 39284 36728 39296
rect 35575 39256 36728 39284
rect 35575 39253 35587 39256
rect 35529 39247 35587 39253
rect 35400 39244 35406 39247
rect 36722 39244 36728 39256
rect 36780 39244 36786 39296
rect 38194 39244 38200 39296
rect 38252 39284 38258 39296
rect 38289 39287 38347 39293
rect 38289 39284 38301 39287
rect 38252 39256 38301 39284
rect 38252 39244 38258 39256
rect 38289 39253 38301 39256
rect 38335 39253 38347 39287
rect 38580 39284 38608 39324
rect 40604 39324 42340 39352
rect 40604 39284 40632 39324
rect 42334 39312 42340 39324
rect 42392 39312 42398 39364
rect 38580 39256 40632 39284
rect 38289 39247 38347 39253
rect 40678 39244 40684 39296
rect 40736 39284 40742 39296
rect 41325 39287 41383 39293
rect 41325 39284 41337 39287
rect 40736 39256 41337 39284
rect 40736 39244 40742 39256
rect 41325 39253 41337 39256
rect 41371 39253 41383 39287
rect 42444 39284 42472 39392
rect 42610 39380 42616 39392
rect 42668 39380 42674 39432
rect 42794 39420 42800 39432
rect 42755 39392 42800 39420
rect 42794 39380 42800 39392
rect 42852 39380 42858 39432
rect 43625 39423 43683 39429
rect 43625 39389 43637 39423
rect 43671 39420 43683 39423
rect 43806 39420 43812 39432
rect 43671 39392 43812 39420
rect 43671 39389 43683 39392
rect 43625 39383 43683 39389
rect 43806 39380 43812 39392
rect 43864 39380 43870 39432
rect 45094 39380 45100 39432
rect 45152 39420 45158 39432
rect 45388 39429 45416 39516
rect 46658 39448 46664 39500
rect 46716 39488 46722 39500
rect 46753 39491 46811 39497
rect 46753 39488 46765 39491
rect 46716 39460 46765 39488
rect 46716 39448 46722 39460
rect 46753 39457 46765 39460
rect 46799 39457 46811 39491
rect 46753 39451 46811 39457
rect 45281 39423 45339 39429
rect 45281 39420 45293 39423
rect 45152 39392 45293 39420
rect 45152 39380 45158 39392
rect 45281 39389 45293 39392
rect 45327 39389 45339 39423
rect 45281 39383 45339 39389
rect 45370 39423 45428 39429
rect 45370 39389 45382 39423
rect 45416 39389 45428 39423
rect 45370 39383 45428 39389
rect 45465 39417 45523 39423
rect 45646 39420 45652 39432
rect 45465 39383 45477 39417
rect 45511 39383 45523 39417
rect 45607 39392 45652 39420
rect 45465 39377 45523 39383
rect 45646 39380 45652 39392
rect 45704 39380 45710 39432
rect 46106 39420 46112 39432
rect 46019 39392 46112 39420
rect 46106 39380 46112 39392
rect 46164 39380 46170 39432
rect 46842 39380 46848 39432
rect 46900 39420 46906 39432
rect 47009 39423 47067 39429
rect 47009 39420 47021 39423
rect 46900 39392 47021 39420
rect 46900 39380 46906 39392
rect 47009 39389 47021 39392
rect 47055 39389 47067 39423
rect 48774 39420 48780 39432
rect 48735 39392 48780 39420
rect 47009 39383 47067 39389
rect 48774 39380 48780 39392
rect 48832 39380 48838 39432
rect 42518 39312 42524 39364
rect 42576 39352 42582 39364
rect 42576 39324 45140 39352
rect 42576 39312 42582 39324
rect 43254 39284 43260 39296
rect 42444 39256 43260 39284
rect 41325 39247 41383 39253
rect 43254 39244 43260 39256
rect 43312 39244 43318 39296
rect 43438 39284 43444 39296
rect 43399 39256 43444 39284
rect 43438 39244 43444 39256
rect 43496 39244 43502 39296
rect 44910 39244 44916 39296
rect 44968 39284 44974 39296
rect 45005 39287 45063 39293
rect 45005 39284 45017 39287
rect 44968 39256 45017 39284
rect 44968 39244 44974 39256
rect 45005 39253 45017 39256
rect 45051 39253 45063 39287
rect 45112 39284 45140 39324
rect 45480 39284 45508 39377
rect 46124 39352 46152 39380
rect 48792 39352 48820 39380
rect 46124 39324 48820 39352
rect 45112 39256 45508 39284
rect 45005 39247 45063 39253
rect 46014 39244 46020 39296
rect 46072 39284 46078 39296
rect 46201 39287 46259 39293
rect 46201 39284 46213 39287
rect 46072 39256 46213 39284
rect 46072 39244 46078 39256
rect 46201 39253 46213 39256
rect 46247 39253 46259 39287
rect 46201 39247 46259 39253
rect 48869 39287 48927 39293
rect 48869 39253 48881 39287
rect 48915 39284 48927 39287
rect 48958 39284 48964 39296
rect 48915 39256 48964 39284
rect 48915 39253 48927 39256
rect 48869 39247 48927 39253
rect 48958 39244 48964 39256
rect 49016 39244 49022 39296
rect 1104 39194 68816 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 68816 39194
rect 1104 39120 68816 39142
rect 1854 39080 1860 39092
rect 1815 39052 1860 39080
rect 1854 39040 1860 39052
rect 1912 39040 1918 39092
rect 19426 39040 19432 39092
rect 19484 39080 19490 39092
rect 19705 39083 19763 39089
rect 19705 39080 19717 39083
rect 19484 39052 19717 39080
rect 19484 39040 19490 39052
rect 19705 39049 19717 39052
rect 19751 39049 19763 39083
rect 22554 39080 22560 39092
rect 22515 39052 22560 39080
rect 19705 39043 19763 39049
rect 22554 39040 22560 39052
rect 22612 39040 22618 39092
rect 23106 39080 23112 39092
rect 22756 39052 23112 39080
rect 1765 38947 1823 38953
rect 1765 38913 1777 38947
rect 1811 38944 1823 38947
rect 3142 38944 3148 38956
rect 1811 38916 3148 38944
rect 1811 38913 1823 38916
rect 1765 38907 1823 38913
rect 3142 38904 3148 38916
rect 3200 38904 3206 38956
rect 19613 38947 19671 38953
rect 19613 38913 19625 38947
rect 19659 38944 19671 38947
rect 19978 38944 19984 38956
rect 19659 38916 19984 38944
rect 19659 38913 19671 38916
rect 19613 38907 19671 38913
rect 19978 38904 19984 38916
rect 20036 38904 20042 38956
rect 20898 38944 20904 38956
rect 20859 38916 20904 38944
rect 20898 38904 20904 38916
rect 20956 38904 20962 38956
rect 20993 38947 21051 38953
rect 20993 38913 21005 38947
rect 21039 38913 21051 38947
rect 20993 38907 21051 38913
rect 21008 38876 21036 38907
rect 21082 38904 21088 38956
rect 21140 38944 21146 38956
rect 21269 38947 21327 38953
rect 21140 38916 21185 38944
rect 21140 38904 21146 38916
rect 21269 38913 21281 38947
rect 21315 38944 21327 38947
rect 22756 38944 22784 39052
rect 23106 39040 23112 39052
rect 23164 39040 23170 39092
rect 26234 39040 26240 39092
rect 26292 39080 26298 39092
rect 27338 39080 27344 39092
rect 26292 39052 27344 39080
rect 26292 39040 26298 39052
rect 27338 39040 27344 39052
rect 27396 39040 27402 39092
rect 28166 39040 28172 39092
rect 28224 39080 28230 39092
rect 28445 39083 28503 39089
rect 28445 39080 28457 39083
rect 28224 39052 28457 39080
rect 28224 39040 28230 39052
rect 28445 39049 28457 39052
rect 28491 39049 28503 39083
rect 31018 39080 31024 39092
rect 30979 39052 31024 39080
rect 28445 39043 28503 39049
rect 22848 38984 23796 39012
rect 22848 38953 22876 38984
rect 23768 38956 23796 38984
rect 25222 38972 25228 39024
rect 25280 39012 25286 39024
rect 26421 39015 26479 39021
rect 26421 39012 26433 39015
rect 25280 38984 26433 39012
rect 25280 38972 25286 38984
rect 26421 38981 26433 38984
rect 26467 39012 26479 39015
rect 28460 39012 28488 39043
rect 31018 39040 31024 39052
rect 31076 39040 31082 39092
rect 35250 39080 35256 39092
rect 35211 39052 35256 39080
rect 35250 39040 35256 39052
rect 35308 39040 35314 39092
rect 38470 39040 38476 39092
rect 38528 39080 38534 39092
rect 39301 39083 39359 39089
rect 39301 39080 39313 39083
rect 38528 39052 39313 39080
rect 38528 39040 38534 39052
rect 39301 39049 39313 39052
rect 39347 39049 39359 39083
rect 40494 39080 40500 39092
rect 40455 39052 40500 39080
rect 39301 39043 39359 39049
rect 40494 39040 40500 39052
rect 40552 39040 40558 39092
rect 42429 39083 42487 39089
rect 42429 39049 42441 39083
rect 42475 39080 42487 39083
rect 42518 39080 42524 39092
rect 42475 39052 42524 39080
rect 42475 39049 42487 39052
rect 42429 39043 42487 39049
rect 42518 39040 42524 39052
rect 42576 39040 42582 39092
rect 43806 39080 43812 39092
rect 43767 39052 43812 39080
rect 43806 39040 43812 39052
rect 43864 39040 43870 39092
rect 45094 39040 45100 39092
rect 45152 39080 45158 39092
rect 45830 39080 45836 39092
rect 45152 39052 45836 39080
rect 45152 39040 45158 39052
rect 45830 39040 45836 39052
rect 45888 39080 45894 39092
rect 46017 39083 46075 39089
rect 46017 39080 46029 39083
rect 45888 39052 46029 39080
rect 45888 39040 45894 39052
rect 46017 39049 46029 39052
rect 46063 39049 46075 39083
rect 46017 39043 46075 39049
rect 39850 39012 39856 39024
rect 26467 38984 28120 39012
rect 28460 38984 33548 39012
rect 26467 38981 26479 38984
rect 26421 38975 26479 38981
rect 21315 38916 22784 38944
rect 22833 38947 22891 38953
rect 21315 38913 21327 38916
rect 21269 38907 21327 38913
rect 22833 38913 22845 38947
rect 22879 38913 22891 38947
rect 22833 38907 22891 38913
rect 22925 38947 22983 38953
rect 22925 38913 22937 38947
rect 22971 38913 22983 38947
rect 22925 38907 22983 38913
rect 22738 38876 22744 38888
rect 21008 38848 22744 38876
rect 22738 38836 22744 38848
rect 22796 38876 22802 38888
rect 22940 38876 22968 38907
rect 23014 38904 23020 38956
rect 23072 38944 23078 38956
rect 23201 38947 23259 38953
rect 23072 38916 23117 38944
rect 23072 38904 23078 38916
rect 23201 38913 23213 38947
rect 23247 38913 23259 38947
rect 23201 38907 23259 38913
rect 22796 38848 22968 38876
rect 22796 38836 22802 38848
rect 23106 38836 23112 38888
rect 23164 38876 23170 38888
rect 23216 38876 23244 38907
rect 23750 38904 23756 38956
rect 23808 38944 23814 38956
rect 23845 38947 23903 38953
rect 23845 38944 23857 38947
rect 23808 38916 23857 38944
rect 23808 38904 23814 38916
rect 23845 38913 23857 38916
rect 23891 38913 23903 38947
rect 26234 38944 26240 38956
rect 26195 38916 26240 38944
rect 23845 38907 23903 38913
rect 26234 38904 26240 38916
rect 26292 38904 26298 38956
rect 27062 38944 27068 38956
rect 27023 38916 27068 38944
rect 27062 38904 27068 38916
rect 27120 38904 27126 38956
rect 27332 38947 27390 38953
rect 27332 38913 27344 38947
rect 27378 38944 27390 38947
rect 27706 38944 27712 38956
rect 27378 38916 27712 38944
rect 27378 38913 27390 38916
rect 27332 38907 27390 38913
rect 27706 38904 27712 38916
rect 27764 38904 27770 38956
rect 24026 38876 24032 38888
rect 23164 38848 23244 38876
rect 23987 38848 24032 38876
rect 23164 38836 23170 38848
rect 24026 38836 24032 38848
rect 24084 38836 24090 38888
rect 25590 38876 25596 38888
rect 25551 38848 25596 38876
rect 25590 38836 25596 38848
rect 25648 38836 25654 38888
rect 28092 38876 28120 38984
rect 30834 38904 30840 38956
rect 30892 38944 30898 38956
rect 30929 38947 30987 38953
rect 30929 38944 30941 38947
rect 30892 38916 30941 38944
rect 30892 38904 30898 38916
rect 30929 38913 30941 38916
rect 30975 38913 30987 38947
rect 32306 38944 32312 38956
rect 30929 38907 30987 38913
rect 31726 38916 32312 38944
rect 31726 38876 31754 38916
rect 32306 38904 32312 38916
rect 32364 38904 32370 38956
rect 33410 38944 33416 38956
rect 33371 38916 33416 38944
rect 33410 38904 33416 38916
rect 33468 38904 33474 38956
rect 33520 38944 33548 38984
rect 37936 38984 39856 39012
rect 35802 38944 35808 38956
rect 33520 38916 33732 38944
rect 35763 38916 35808 38944
rect 28092 38848 31754 38876
rect 32125 38879 32183 38885
rect 32125 38845 32137 38879
rect 32171 38876 32183 38879
rect 33594 38876 33600 38888
rect 32171 38848 32904 38876
rect 33555 38848 33600 38876
rect 32171 38845 32183 38848
rect 32125 38839 32183 38845
rect 32876 38752 32904 38848
rect 33594 38836 33600 38848
rect 33652 38836 33658 38888
rect 33704 38876 33732 38916
rect 35802 38904 35808 38916
rect 35860 38904 35866 38956
rect 36722 38944 36728 38956
rect 36683 38916 36728 38944
rect 36722 38904 36728 38916
rect 36780 38904 36786 38956
rect 37936 38953 37964 38984
rect 39850 38972 39856 38984
rect 39908 38972 39914 39024
rect 41046 38972 41052 39024
rect 41104 39012 41110 39024
rect 41601 39015 41659 39021
rect 41601 39012 41613 39015
rect 41104 38984 41613 39012
rect 41104 38972 41110 38984
rect 41601 38981 41613 38984
rect 41647 38981 41659 39015
rect 41601 38975 41659 38981
rect 43254 38972 43260 39024
rect 43312 39012 43318 39024
rect 43714 39012 43720 39024
rect 43312 38984 43720 39012
rect 43312 38972 43318 38984
rect 38194 38953 38200 38956
rect 37921 38947 37979 38953
rect 37921 38913 37933 38947
rect 37967 38913 37979 38947
rect 38188 38944 38200 38953
rect 38155 38916 38200 38944
rect 37921 38907 37979 38913
rect 38188 38907 38200 38916
rect 38194 38904 38200 38907
rect 38252 38904 38258 38956
rect 40678 38944 40684 38956
rect 40639 38916 40684 38944
rect 40678 38904 40684 38916
rect 40736 38904 40742 38956
rect 41414 38904 41420 38956
rect 41472 38944 41478 38956
rect 41472 38916 41517 38944
rect 41472 38904 41478 38916
rect 42334 38904 42340 38956
rect 42392 38944 42398 38956
rect 42705 38947 42763 38953
rect 42705 38944 42717 38947
rect 42392 38916 42717 38944
rect 42392 38904 42398 38916
rect 42705 38913 42717 38916
rect 42751 38913 42763 38947
rect 42886 38944 42892 38956
rect 42847 38916 42892 38944
rect 42705 38907 42763 38913
rect 42886 38904 42892 38916
rect 42944 38904 42950 38956
rect 43346 38904 43352 38956
rect 43404 38944 43410 38956
rect 43640 38953 43668 38984
rect 43714 38972 43720 38984
rect 43772 38972 43778 39024
rect 45186 39012 45192 39024
rect 44652 38984 45192 39012
rect 44652 38953 44680 38984
rect 45186 38972 45192 38984
rect 45244 39012 45250 39024
rect 46658 39012 46664 39024
rect 45244 38984 46664 39012
rect 45244 38972 45250 38984
rect 46658 38972 46664 38984
rect 46716 38972 46722 39024
rect 48958 39012 48964 39024
rect 48919 38984 48964 39012
rect 48958 38972 48964 38984
rect 49016 38972 49022 39024
rect 44910 38953 44916 38956
rect 43441 38947 43499 38953
rect 43441 38944 43453 38947
rect 43404 38916 43453 38944
rect 43404 38904 43410 38916
rect 43441 38913 43453 38916
rect 43487 38913 43499 38947
rect 43441 38907 43499 38913
rect 43625 38947 43683 38953
rect 43625 38913 43637 38947
rect 43671 38913 43683 38947
rect 43625 38907 43683 38913
rect 44637 38947 44695 38953
rect 44637 38913 44649 38947
rect 44683 38913 44695 38947
rect 44904 38944 44916 38953
rect 44871 38916 44916 38944
rect 44637 38907 44695 38913
rect 44904 38907 44916 38916
rect 34333 38879 34391 38885
rect 34333 38876 34345 38879
rect 33704 38848 34345 38876
rect 34333 38845 34345 38848
rect 34379 38845 34391 38879
rect 34333 38839 34391 38845
rect 34422 38836 34428 38888
rect 34480 38885 34486 38888
rect 34480 38879 34508 38885
rect 34496 38845 34508 38879
rect 34480 38839 34508 38845
rect 34609 38879 34667 38885
rect 34609 38845 34621 38879
rect 34655 38876 34667 38879
rect 34790 38876 34796 38888
rect 34655 38848 34796 38876
rect 34655 38845 34667 38848
rect 34609 38839 34667 38845
rect 34480 38836 34486 38839
rect 34790 38836 34796 38848
rect 34848 38876 34854 38888
rect 35342 38876 35348 38888
rect 34848 38848 35348 38876
rect 34848 38836 34854 38848
rect 35342 38836 35348 38848
rect 35400 38836 35406 38888
rect 41785 38879 41843 38885
rect 41785 38845 41797 38879
rect 41831 38876 41843 38879
rect 42613 38879 42671 38885
rect 42613 38876 42625 38879
rect 41831 38848 42625 38876
rect 41831 38845 41843 38848
rect 41785 38839 41843 38845
rect 42613 38845 42625 38848
rect 42659 38845 42671 38879
rect 42794 38876 42800 38888
rect 42755 38848 42800 38876
rect 42613 38839 42671 38845
rect 42794 38836 42800 38848
rect 42852 38836 42858 38888
rect 33870 38768 33876 38820
rect 33928 38808 33934 38820
rect 34054 38808 34060 38820
rect 33928 38780 34060 38808
rect 33928 38768 33934 38780
rect 34054 38768 34060 38780
rect 34112 38768 34118 38820
rect 42702 38768 42708 38820
rect 42760 38808 42766 38820
rect 42904 38808 42932 38904
rect 43456 38876 43484 38907
rect 44910 38904 44916 38907
rect 44968 38904 44974 38956
rect 48038 38904 48044 38956
rect 48096 38944 48102 38956
rect 48777 38947 48835 38953
rect 48777 38944 48789 38947
rect 48096 38916 48789 38944
rect 48096 38904 48102 38916
rect 48777 38913 48789 38916
rect 48823 38913 48835 38947
rect 48777 38907 48835 38913
rect 44082 38876 44088 38888
rect 43456 38848 44088 38876
rect 44082 38836 44088 38848
rect 44140 38836 44146 38888
rect 50614 38876 50620 38888
rect 50575 38848 50620 38876
rect 50614 38836 50620 38848
rect 50672 38836 50678 38888
rect 42760 38780 42932 38808
rect 42760 38768 42766 38780
rect 20625 38743 20683 38749
rect 20625 38709 20637 38743
rect 20671 38740 20683 38743
rect 21174 38740 21180 38752
rect 20671 38712 21180 38740
rect 20671 38709 20683 38712
rect 20625 38703 20683 38709
rect 21174 38700 21180 38712
rect 21232 38700 21238 38752
rect 32306 38700 32312 38752
rect 32364 38740 32370 38752
rect 32493 38743 32551 38749
rect 32493 38740 32505 38743
rect 32364 38712 32505 38740
rect 32364 38700 32370 38712
rect 32493 38709 32505 38712
rect 32539 38709 32551 38743
rect 32493 38703 32551 38709
rect 32858 38700 32864 38752
rect 32916 38740 32922 38752
rect 34422 38740 34428 38752
rect 32916 38712 34428 38740
rect 32916 38700 32922 38712
rect 34422 38700 34428 38712
rect 34480 38700 34486 38752
rect 35986 38740 35992 38752
rect 35947 38712 35992 38740
rect 35986 38700 35992 38712
rect 36044 38700 36050 38752
rect 36538 38740 36544 38752
rect 36499 38712 36544 38740
rect 36538 38700 36544 38712
rect 36596 38700 36602 38752
rect 1104 38650 68816 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 65654 38650
rect 65706 38598 65718 38650
rect 65770 38598 65782 38650
rect 65834 38598 65846 38650
rect 65898 38598 65910 38650
rect 65962 38598 68816 38650
rect 1104 38576 68816 38598
rect 3234 38496 3240 38548
rect 3292 38536 3298 38548
rect 20714 38536 20720 38548
rect 3292 38508 20720 38536
rect 3292 38496 3298 38508
rect 20714 38496 20720 38508
rect 20772 38496 20778 38548
rect 23661 38539 23719 38545
rect 23661 38505 23673 38539
rect 23707 38536 23719 38539
rect 24026 38536 24032 38548
rect 23707 38508 24032 38536
rect 23707 38505 23719 38508
rect 23661 38499 23719 38505
rect 24026 38496 24032 38508
rect 24084 38496 24090 38548
rect 27706 38536 27712 38548
rect 27667 38508 27712 38536
rect 27706 38496 27712 38508
rect 27764 38496 27770 38548
rect 32769 38539 32827 38545
rect 32769 38505 32781 38539
rect 32815 38536 32827 38539
rect 32858 38536 32864 38548
rect 32815 38508 32864 38536
rect 32815 38505 32827 38508
rect 32769 38499 32827 38505
rect 32858 38496 32864 38508
rect 32916 38496 32922 38548
rect 35434 38496 35440 38548
rect 35492 38536 35498 38548
rect 36909 38539 36967 38545
rect 36909 38536 36921 38539
rect 35492 38508 36921 38536
rect 35492 38496 35498 38508
rect 36909 38505 36921 38508
rect 36955 38505 36967 38539
rect 36909 38499 36967 38505
rect 39850 38496 39856 38548
rect 39908 38536 39914 38548
rect 41601 38539 41659 38545
rect 41601 38536 41613 38539
rect 39908 38508 41613 38536
rect 39908 38496 39914 38508
rect 41601 38505 41613 38508
rect 41647 38536 41659 38539
rect 45186 38536 45192 38548
rect 41647 38508 45192 38536
rect 41647 38505 41659 38508
rect 41601 38499 41659 38505
rect 45186 38496 45192 38508
rect 45244 38496 45250 38548
rect 44082 38428 44088 38480
rect 44140 38468 44146 38480
rect 44269 38471 44327 38477
rect 44269 38468 44281 38471
rect 44140 38440 44281 38468
rect 44140 38428 44146 38440
rect 44269 38437 44281 38440
rect 44315 38437 44327 38471
rect 44269 38431 44327 38437
rect 37366 38400 37372 38412
rect 37327 38372 37372 38400
rect 37366 38360 37372 38372
rect 37424 38360 37430 38412
rect 45830 38400 45836 38412
rect 45791 38372 45836 38400
rect 45830 38360 45836 38372
rect 45888 38360 45894 38412
rect 46014 38400 46020 38412
rect 45975 38372 46020 38400
rect 46014 38360 46020 38372
rect 46072 38360 46078 38412
rect 19797 38335 19855 38341
rect 19797 38301 19809 38335
rect 19843 38332 19855 38335
rect 19978 38332 19984 38344
rect 19843 38304 19984 38332
rect 19843 38301 19855 38304
rect 19797 38295 19855 38301
rect 19978 38292 19984 38304
rect 20036 38292 20042 38344
rect 20901 38335 20959 38341
rect 20901 38301 20913 38335
rect 20947 38332 20959 38335
rect 22370 38332 22376 38344
rect 20947 38304 22376 38332
rect 20947 38301 20959 38304
rect 20901 38295 20959 38301
rect 22370 38292 22376 38304
rect 22428 38292 22434 38344
rect 23382 38292 23388 38344
rect 23440 38332 23446 38344
rect 23569 38335 23627 38341
rect 23569 38332 23581 38335
rect 23440 38304 23581 38332
rect 23440 38292 23446 38304
rect 23569 38301 23581 38304
rect 23615 38301 23627 38335
rect 24394 38332 24400 38344
rect 24355 38304 24400 38332
rect 23569 38295 23627 38301
rect 24394 38292 24400 38304
rect 24452 38292 24458 38344
rect 27890 38332 27896 38344
rect 27851 38304 27896 38332
rect 27890 38292 27896 38304
rect 27948 38292 27954 38344
rect 29825 38335 29883 38341
rect 29825 38301 29837 38335
rect 29871 38332 29883 38335
rect 30190 38332 30196 38344
rect 29871 38304 30196 38332
rect 29871 38301 29883 38304
rect 29825 38295 29883 38301
rect 30190 38292 30196 38304
rect 30248 38292 30254 38344
rect 30834 38332 30840 38344
rect 30795 38304 30840 38332
rect 30834 38292 30840 38304
rect 30892 38292 30898 38344
rect 30929 38335 30987 38341
rect 30929 38301 30941 38335
rect 30975 38332 30987 38335
rect 31389 38335 31447 38341
rect 31389 38332 31401 38335
rect 30975 38304 31401 38332
rect 30975 38301 30987 38304
rect 30929 38295 30987 38301
rect 31389 38301 31401 38304
rect 31435 38301 31447 38335
rect 31389 38295 31447 38301
rect 34977 38335 35035 38341
rect 34977 38301 34989 38335
rect 35023 38301 35035 38335
rect 34977 38295 35035 38301
rect 35069 38335 35127 38341
rect 35069 38301 35081 38335
rect 35115 38332 35127 38335
rect 35529 38335 35587 38341
rect 35529 38332 35541 38335
rect 35115 38304 35541 38332
rect 35115 38301 35127 38304
rect 35069 38295 35127 38301
rect 35529 38301 35541 38304
rect 35575 38301 35587 38335
rect 35529 38295 35587 38301
rect 35796 38335 35854 38341
rect 35796 38301 35808 38335
rect 35842 38332 35854 38335
rect 36538 38332 36544 38344
rect 35842 38304 36544 38332
rect 35842 38301 35854 38304
rect 35796 38295 35854 38301
rect 21174 38273 21180 38276
rect 21168 38264 21180 38273
rect 21135 38236 21180 38264
rect 21168 38227 21180 38236
rect 21174 38224 21180 38227
rect 21232 38224 21238 38276
rect 24670 38273 24676 38276
rect 24664 38227 24676 38273
rect 24728 38264 24734 38276
rect 31656 38267 31714 38273
rect 24728 38236 24764 38264
rect 24670 38224 24676 38227
rect 24728 38224 24734 38236
rect 31656 38233 31668 38267
rect 31702 38264 31714 38267
rect 32122 38264 32128 38276
rect 31702 38236 32128 38264
rect 31702 38233 31714 38236
rect 31656 38227 31714 38233
rect 32122 38224 32128 38236
rect 32180 38224 32186 38276
rect 33778 38264 33784 38276
rect 33739 38236 33784 38264
rect 33778 38224 33784 38236
rect 33836 38224 33842 38276
rect 33965 38267 34023 38273
rect 33965 38233 33977 38267
rect 34011 38264 34023 38267
rect 34054 38264 34060 38276
rect 34011 38236 34060 38264
rect 34011 38233 34023 38236
rect 33965 38227 34023 38233
rect 34054 38224 34060 38236
rect 34112 38264 34118 38276
rect 34514 38264 34520 38276
rect 34112 38236 34520 38264
rect 34112 38224 34118 38236
rect 34514 38224 34520 38236
rect 34572 38224 34578 38276
rect 34992 38264 35020 38295
rect 36538 38292 36544 38304
rect 36596 38292 36602 38344
rect 37642 38332 37648 38344
rect 37603 38304 37648 38332
rect 37642 38292 37648 38304
rect 37700 38292 37706 38344
rect 38378 38292 38384 38344
rect 38436 38332 38442 38344
rect 40405 38335 40463 38341
rect 40405 38332 40417 38335
rect 38436 38304 40417 38332
rect 38436 38292 38442 38304
rect 40405 38301 40417 38304
rect 40451 38301 40463 38335
rect 40405 38295 40463 38301
rect 40954 38292 40960 38344
rect 41012 38332 41018 38344
rect 42153 38335 42211 38341
rect 42153 38332 42165 38335
rect 41012 38304 42165 38332
rect 41012 38292 41018 38304
rect 42153 38301 42165 38304
rect 42199 38301 42211 38335
rect 42153 38295 42211 38301
rect 42429 38335 42487 38341
rect 42429 38301 42441 38335
rect 42475 38332 42487 38335
rect 42889 38335 42947 38341
rect 42889 38332 42901 38335
rect 42475 38304 42901 38332
rect 42475 38301 42487 38304
rect 42429 38295 42487 38301
rect 42889 38301 42901 38304
rect 42935 38301 42947 38335
rect 42889 38295 42947 38301
rect 43156 38335 43214 38341
rect 43156 38301 43168 38335
rect 43202 38332 43214 38335
rect 43438 38332 43444 38344
rect 43202 38304 43444 38332
rect 43202 38301 43214 38304
rect 43156 38295 43214 38301
rect 43438 38292 43444 38304
rect 43496 38292 43502 38344
rect 50157 38335 50215 38341
rect 50157 38332 50169 38335
rect 47504 38304 50169 38332
rect 35986 38264 35992 38276
rect 34992 38236 35992 38264
rect 35986 38224 35992 38236
rect 36044 38224 36050 38276
rect 40586 38264 40592 38276
rect 40547 38236 40592 38264
rect 40586 38224 40592 38236
rect 40644 38264 40650 38276
rect 41509 38267 41567 38273
rect 41509 38264 41521 38267
rect 40644 38236 41521 38264
rect 40644 38224 40650 38236
rect 41509 38233 41521 38236
rect 41555 38233 41567 38267
rect 47504 38264 47532 38304
rect 50157 38301 50169 38304
rect 50203 38332 50215 38335
rect 66806 38332 66812 38344
rect 50203 38304 66812 38332
rect 50203 38301 50215 38304
rect 50157 38295 50215 38301
rect 66806 38292 66812 38304
rect 66864 38292 66870 38344
rect 41509 38227 41567 38233
rect 44192 38236 47532 38264
rect 19889 38199 19947 38205
rect 19889 38165 19901 38199
rect 19935 38196 19947 38199
rect 19978 38196 19984 38208
rect 19935 38168 19984 38196
rect 19935 38165 19947 38168
rect 19889 38159 19947 38165
rect 19978 38156 19984 38168
rect 20036 38156 20042 38208
rect 20898 38156 20904 38208
rect 20956 38196 20962 38208
rect 22281 38199 22339 38205
rect 22281 38196 22293 38199
rect 20956 38168 22293 38196
rect 20956 38156 20962 38168
rect 22281 38165 22293 38168
rect 22327 38165 22339 38199
rect 22281 38159 22339 38165
rect 25777 38199 25835 38205
rect 25777 38165 25789 38199
rect 25823 38196 25835 38199
rect 27246 38196 27252 38208
rect 25823 38168 27252 38196
rect 25823 38165 25835 38168
rect 25777 38159 25835 38165
rect 27246 38156 27252 38168
rect 27304 38156 27310 38208
rect 29638 38196 29644 38208
rect 29599 38168 29644 38196
rect 29638 38156 29644 38168
rect 29696 38156 29702 38208
rect 32214 38156 32220 38208
rect 32272 38196 32278 38208
rect 44192 38196 44220 38236
rect 47578 38224 47584 38276
rect 47636 38264 47642 38276
rect 47673 38267 47731 38273
rect 47673 38264 47685 38267
rect 47636 38236 47685 38264
rect 47636 38224 47642 38236
rect 47673 38233 47685 38236
rect 47719 38233 47731 38267
rect 47673 38227 47731 38233
rect 32272 38168 44220 38196
rect 32272 38156 32278 38168
rect 50062 38156 50068 38208
rect 50120 38196 50126 38208
rect 50249 38199 50307 38205
rect 50249 38196 50261 38199
rect 50120 38168 50261 38196
rect 50120 38156 50126 38168
rect 50249 38165 50261 38168
rect 50295 38165 50307 38199
rect 50249 38159 50307 38165
rect 66622 38156 66628 38208
rect 66680 38196 66686 38208
rect 66806 38196 66812 38208
rect 66680 38168 66812 38196
rect 66680 38156 66686 38168
rect 66806 38156 66812 38168
rect 66864 38156 66870 38208
rect 1104 38106 68816 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 68816 38106
rect 1104 38032 68816 38054
rect 20898 37992 20904 38004
rect 19444 37964 20904 37992
rect 19444 37865 19472 37964
rect 20898 37952 20904 37964
rect 20956 37952 20962 38004
rect 24394 37952 24400 38004
rect 24452 37992 24458 38004
rect 25317 37995 25375 38001
rect 25317 37992 25329 37995
rect 24452 37964 25329 37992
rect 24452 37952 24458 37964
rect 25317 37961 25329 37964
rect 25363 37961 25375 37995
rect 32122 37992 32128 38004
rect 32083 37964 32128 37992
rect 25317 37955 25375 37961
rect 32122 37952 32128 37964
rect 32180 37952 32186 38004
rect 38562 37952 38568 38004
rect 38620 37992 38626 38004
rect 40862 37992 40868 38004
rect 38620 37964 40868 37992
rect 38620 37952 38626 37964
rect 40862 37952 40868 37964
rect 40920 37992 40926 38004
rect 40920 37964 41414 37992
rect 40920 37952 40926 37964
rect 19613 37927 19671 37933
rect 19613 37893 19625 37927
rect 19659 37924 19671 37927
rect 19978 37924 19984 37936
rect 19659 37896 19984 37924
rect 19659 37893 19671 37896
rect 19613 37887 19671 37893
rect 19978 37884 19984 37896
rect 20036 37884 20042 37936
rect 27154 37924 27160 37936
rect 27115 37896 27160 37924
rect 27154 37884 27160 37896
rect 27212 37884 27218 37936
rect 27373 37927 27431 37933
rect 27373 37893 27385 37927
rect 27419 37924 27431 37927
rect 28810 37924 28816 37936
rect 27419 37896 28816 37924
rect 27419 37893 27431 37896
rect 27373 37887 27431 37893
rect 28810 37884 28816 37896
rect 28868 37884 28874 37936
rect 29638 37933 29644 37936
rect 29632 37924 29644 37933
rect 29599 37896 29644 37924
rect 29632 37887 29644 37896
rect 29638 37884 29644 37887
rect 29696 37884 29702 37936
rect 37458 37884 37464 37936
rect 37516 37924 37522 37936
rect 37737 37927 37795 37933
rect 37737 37924 37749 37927
rect 37516 37896 37749 37924
rect 37516 37884 37522 37896
rect 37737 37893 37749 37896
rect 37783 37893 37795 37927
rect 38746 37924 38752 37936
rect 38707 37896 38752 37924
rect 37737 37887 37795 37893
rect 38746 37884 38752 37896
rect 38804 37884 38810 37936
rect 39942 37884 39948 37936
rect 40000 37924 40006 37936
rect 40098 37927 40156 37933
rect 40098 37924 40110 37927
rect 40000 37896 40110 37924
rect 40000 37884 40006 37896
rect 40098 37893 40110 37896
rect 40144 37893 40156 37927
rect 40098 37887 40156 37893
rect 19429 37859 19487 37865
rect 19429 37825 19441 37859
rect 19475 37825 19487 37859
rect 23290 37856 23296 37868
rect 23251 37828 23296 37856
rect 19429 37819 19487 37825
rect 23290 37816 23296 37828
rect 23348 37816 23354 37868
rect 25317 37859 25375 37865
rect 25317 37825 25329 37859
rect 25363 37856 25375 37859
rect 25774 37856 25780 37868
rect 25363 37828 25780 37856
rect 25363 37825 25375 37828
rect 25317 37819 25375 37825
rect 25774 37816 25780 37828
rect 25832 37816 25838 37868
rect 26050 37856 26056 37868
rect 25963 37828 26056 37856
rect 26050 37816 26056 37828
rect 26108 37856 26114 37868
rect 26418 37856 26424 37868
rect 26108 37828 26424 37856
rect 26108 37816 26114 37828
rect 26418 37816 26424 37828
rect 26476 37816 26482 37868
rect 29362 37856 29368 37868
rect 29323 37828 29368 37856
rect 29362 37816 29368 37828
rect 29420 37816 29426 37868
rect 32306 37856 32312 37868
rect 32267 37828 32312 37856
rect 32306 37816 32312 37828
rect 32364 37816 32370 37868
rect 32674 37816 32680 37868
rect 32732 37856 32738 37868
rect 32861 37859 32919 37865
rect 32861 37856 32873 37859
rect 32732 37828 32873 37856
rect 32732 37816 32738 37828
rect 32861 37825 32873 37828
rect 32907 37856 32919 37859
rect 33318 37856 33324 37868
rect 32907 37828 33324 37856
rect 32907 37825 32919 37828
rect 32861 37819 32919 37825
rect 33318 37816 33324 37828
rect 33376 37816 33382 37868
rect 35529 37859 35587 37865
rect 35529 37825 35541 37859
rect 35575 37856 35587 37859
rect 35802 37856 35808 37868
rect 35575 37828 35808 37856
rect 35575 37825 35587 37828
rect 35529 37819 35587 37825
rect 35802 37816 35808 37828
rect 35860 37816 35866 37868
rect 37550 37856 37556 37868
rect 37511 37828 37556 37856
rect 37550 37816 37556 37828
rect 37608 37816 37614 37868
rect 39002 37856 39008 37868
rect 38963 37828 39008 37856
rect 39002 37816 39008 37828
rect 39060 37816 39066 37868
rect 39117 37859 39175 37865
rect 39117 37825 39129 37859
rect 39163 37825 39175 37859
rect 39117 37819 39175 37825
rect 39209 37862 39267 37868
rect 39209 37828 39221 37862
rect 39255 37828 39267 37862
rect 39209 37822 39267 37828
rect 39393 37859 39451 37865
rect 39393 37825 39405 37859
rect 39439 37856 39451 37859
rect 39482 37856 39488 37868
rect 39439 37828 39488 37856
rect 39439 37825 39451 37828
rect 19889 37791 19947 37797
rect 19889 37757 19901 37791
rect 19935 37757 19947 37791
rect 24210 37788 24216 37800
rect 24171 37760 24216 37788
rect 19889 37751 19947 37757
rect 14 37680 20 37732
rect 72 37720 78 37732
rect 19904 37720 19932 37751
rect 24210 37748 24216 37760
rect 24268 37788 24274 37800
rect 26142 37788 26148 37800
rect 24268 37760 26148 37788
rect 24268 37748 24274 37760
rect 26142 37748 26148 37760
rect 26200 37748 26206 37800
rect 33137 37791 33195 37797
rect 33137 37757 33149 37791
rect 33183 37788 33195 37791
rect 33226 37788 33232 37800
rect 33183 37760 33232 37788
rect 33183 37757 33195 37760
rect 33137 37751 33195 37757
rect 33226 37748 33232 37760
rect 33284 37748 33290 37800
rect 34698 37748 34704 37800
rect 34756 37788 34762 37800
rect 35713 37791 35771 37797
rect 35713 37788 35725 37791
rect 34756 37760 35725 37788
rect 34756 37748 34762 37760
rect 35713 37757 35725 37760
rect 35759 37757 35771 37791
rect 39123 37788 39151 37819
rect 39224 37788 39252 37822
rect 39393 37819 39451 37825
rect 39482 37816 39488 37828
rect 39540 37816 39546 37868
rect 39850 37856 39856 37868
rect 39811 37828 39856 37856
rect 39850 37816 39856 37828
rect 39908 37816 39914 37868
rect 41386 37856 41414 37964
rect 44358 37924 44364 37936
rect 44319 37896 44364 37924
rect 44358 37884 44364 37896
rect 44416 37884 44422 37936
rect 47302 37884 47308 37936
rect 47360 37924 47366 37936
rect 48038 37924 48044 37936
rect 47360 37896 48044 37924
rect 47360 37884 47366 37896
rect 48038 37884 48044 37896
rect 48096 37884 48102 37936
rect 50062 37924 50068 37936
rect 50023 37896 50068 37924
rect 50062 37884 50068 37896
rect 50120 37884 50126 37936
rect 42429 37859 42487 37865
rect 42429 37856 42441 37859
rect 41386 37828 42441 37856
rect 42429 37825 42441 37828
rect 42475 37825 42487 37859
rect 42702 37856 42708 37868
rect 42663 37828 42708 37856
rect 42429 37819 42487 37825
rect 42702 37816 42708 37828
rect 42760 37816 42766 37868
rect 45002 37856 45008 37868
rect 44963 37828 45008 37856
rect 45002 37816 45008 37828
rect 45060 37816 45066 37868
rect 39298 37788 39304 37800
rect 39123 37760 39160 37788
rect 39224 37760 39304 37788
rect 35713 37751 35771 37757
rect 35434 37720 35440 37732
rect 72 37692 19932 37720
rect 30300 37692 35440 37720
rect 72 37680 78 37692
rect 25314 37612 25320 37664
rect 25372 37652 25378 37664
rect 25869 37655 25927 37661
rect 25869 37652 25881 37655
rect 25372 37624 25881 37652
rect 25372 37612 25378 37624
rect 25869 37621 25881 37624
rect 25915 37621 25927 37655
rect 27338 37652 27344 37664
rect 27299 37624 27344 37652
rect 25869 37615 25927 37621
rect 27338 37612 27344 37624
rect 27396 37612 27402 37664
rect 27522 37652 27528 37664
rect 27483 37624 27528 37652
rect 27522 37612 27528 37624
rect 27580 37612 27586 37664
rect 30006 37612 30012 37664
rect 30064 37652 30070 37664
rect 30300 37652 30328 37692
rect 35434 37680 35440 37692
rect 35492 37680 35498 37732
rect 37921 37723 37979 37729
rect 37921 37689 37933 37723
rect 37967 37720 37979 37723
rect 39022 37720 39028 37732
rect 37967 37692 39028 37720
rect 37967 37689 37979 37692
rect 37921 37683 37979 37689
rect 39022 37680 39028 37692
rect 39080 37680 39086 37732
rect 39132 37720 39160 37760
rect 39298 37748 39304 37760
rect 39356 37748 39362 37800
rect 46566 37748 46572 37800
rect 46624 37788 46630 37800
rect 47581 37791 47639 37797
rect 47581 37788 47593 37791
rect 46624 37760 47593 37788
rect 46624 37748 46630 37760
rect 47581 37757 47593 37760
rect 47627 37757 47639 37791
rect 47762 37788 47768 37800
rect 47723 37760 47768 37788
rect 47581 37751 47639 37757
rect 47762 37748 47768 37760
rect 47820 37748 47826 37800
rect 48038 37788 48044 37800
rect 47999 37760 48044 37788
rect 48038 37748 48044 37760
rect 48096 37748 48102 37800
rect 49881 37791 49939 37797
rect 49881 37757 49893 37791
rect 49927 37757 49939 37791
rect 51718 37788 51724 37800
rect 51679 37760 51724 37788
rect 49881 37751 49939 37757
rect 39850 37720 39856 37732
rect 39132 37692 39856 37720
rect 39850 37680 39856 37692
rect 39908 37680 39914 37732
rect 41233 37723 41291 37729
rect 41233 37689 41245 37723
rect 41279 37720 41291 37723
rect 49896 37720 49924 37751
rect 51718 37748 51724 37760
rect 51776 37748 51782 37800
rect 41279 37692 49924 37720
rect 41279 37689 41291 37692
rect 41233 37683 41291 37689
rect 30064 37624 30328 37652
rect 30064 37612 30070 37624
rect 30374 37612 30380 37664
rect 30432 37652 30438 37664
rect 30745 37655 30803 37661
rect 30745 37652 30757 37655
rect 30432 37624 30757 37652
rect 30432 37612 30438 37624
rect 30745 37621 30757 37624
rect 30791 37621 30803 37655
rect 30745 37615 30803 37621
rect 38930 37612 38936 37664
rect 38988 37652 38994 37664
rect 41248 37652 41276 37683
rect 38988 37624 41276 37652
rect 44453 37655 44511 37661
rect 38988 37612 38994 37624
rect 44453 37621 44465 37655
rect 44499 37652 44511 37655
rect 44910 37652 44916 37664
rect 44499 37624 44916 37652
rect 44499 37621 44511 37624
rect 44453 37615 44511 37621
rect 44910 37612 44916 37624
rect 44968 37612 44974 37664
rect 45189 37655 45247 37661
rect 45189 37621 45201 37655
rect 45235 37652 45247 37655
rect 46842 37652 46848 37664
rect 45235 37624 46848 37652
rect 45235 37621 45247 37624
rect 45189 37615 45247 37621
rect 46842 37612 46848 37624
rect 46900 37612 46906 37664
rect 1104 37562 68816 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 68816 37562
rect 1104 37488 68816 37510
rect 27246 37448 27252 37460
rect 24504 37420 27252 37448
rect 24504 37321 24532 37420
rect 27246 37408 27252 37420
rect 27304 37408 27310 37460
rect 28997 37451 29055 37457
rect 28997 37417 29009 37451
rect 29043 37448 29055 37451
rect 37550 37448 37556 37460
rect 29043 37420 37556 37448
rect 29043 37417 29055 37420
rect 28997 37411 29055 37417
rect 37550 37408 37556 37420
rect 37608 37408 37614 37460
rect 38749 37451 38807 37457
rect 38749 37417 38761 37451
rect 38795 37448 38807 37451
rect 39298 37448 39304 37460
rect 38795 37420 39304 37448
rect 38795 37417 38807 37420
rect 38749 37411 38807 37417
rect 39298 37408 39304 37420
rect 39356 37408 39362 37460
rect 39482 37408 39488 37460
rect 39540 37448 39546 37460
rect 40678 37448 40684 37460
rect 39540 37420 40684 37448
rect 39540 37408 39546 37420
rect 40678 37408 40684 37420
rect 40736 37408 40742 37460
rect 47305 37451 47363 37457
rect 47305 37417 47317 37451
rect 47351 37448 47363 37451
rect 47762 37448 47768 37460
rect 47351 37420 47768 37448
rect 47351 37417 47363 37420
rect 47305 37411 47363 37417
rect 47762 37408 47768 37420
rect 47820 37408 47826 37460
rect 26697 37383 26755 37389
rect 26697 37349 26709 37383
rect 26743 37349 26755 37383
rect 26697 37343 26755 37349
rect 22465 37315 22523 37321
rect 22465 37312 22477 37315
rect 21928 37284 22477 37312
rect 3234 37136 3240 37188
rect 3292 37176 3298 37188
rect 21928 37176 21956 37284
rect 22465 37281 22477 37284
rect 22511 37281 22523 37315
rect 22465 37275 22523 37281
rect 24489 37315 24547 37321
rect 24489 37281 24501 37315
rect 24535 37281 24547 37315
rect 25314 37312 25320 37324
rect 25275 37284 25320 37312
rect 24489 37275 24547 37281
rect 25314 37272 25320 37284
rect 25372 37272 25378 37324
rect 26712 37312 26740 37343
rect 27706 37340 27712 37392
rect 27764 37380 27770 37392
rect 27801 37383 27859 37389
rect 27801 37380 27813 37383
rect 27764 37352 27813 37380
rect 27764 37340 27770 37352
rect 27801 37349 27813 37352
rect 27847 37380 27859 37383
rect 27890 37380 27896 37392
rect 27847 37352 27896 37380
rect 27847 37349 27859 37352
rect 27801 37343 27859 37349
rect 27890 37340 27896 37352
rect 27948 37340 27954 37392
rect 30006 37340 30012 37392
rect 30064 37340 30070 37392
rect 43070 37380 43076 37392
rect 41386 37352 43076 37380
rect 27154 37312 27160 37324
rect 26712 37284 27160 37312
rect 27154 37272 27160 37284
rect 27212 37272 27218 37324
rect 27246 37272 27252 37324
rect 27304 37312 27310 37324
rect 28194 37315 28252 37321
rect 28194 37312 28206 37315
rect 27304 37284 28206 37312
rect 27304 37272 27310 37284
rect 28194 37281 28206 37284
rect 28240 37281 28252 37315
rect 28194 37275 28252 37281
rect 29733 37315 29791 37321
rect 29733 37281 29745 37315
rect 29779 37312 29791 37315
rect 30024 37312 30052 37340
rect 35434 37312 35440 37324
rect 29779 37284 30052 37312
rect 35395 37284 35440 37312
rect 29779 37281 29791 37284
rect 29733 37275 29791 37281
rect 35434 37272 35440 37284
rect 35492 37272 35498 37324
rect 35618 37272 35624 37324
rect 35676 37312 35682 37324
rect 35986 37312 35992 37324
rect 35676 37284 35992 37312
rect 35676 37272 35682 37284
rect 35986 37272 35992 37284
rect 36044 37312 36050 37324
rect 39114 37312 39120 37324
rect 36044 37284 36768 37312
rect 39027 37284 39120 37312
rect 36044 37272 36050 37284
rect 22005 37247 22063 37253
rect 22005 37213 22017 37247
rect 22051 37213 22063 37247
rect 22005 37207 22063 37213
rect 24673 37247 24731 37253
rect 24673 37213 24685 37247
rect 24719 37244 24731 37247
rect 27341 37247 27399 37253
rect 24719 37216 25544 37244
rect 24719 37213 24731 37216
rect 24673 37207 24731 37213
rect 3292 37148 21956 37176
rect 3292 37136 3298 37148
rect 22020 37108 22048 37207
rect 22189 37179 22247 37185
rect 22189 37145 22201 37179
rect 22235 37176 22247 37179
rect 22738 37176 22744 37188
rect 22235 37148 22744 37176
rect 22235 37145 22247 37148
rect 22189 37139 22247 37145
rect 22738 37136 22744 37148
rect 22796 37136 22802 37188
rect 25516 37120 25544 37216
rect 27341 37213 27353 37247
rect 27387 37213 27399 37247
rect 27341 37207 27399 37213
rect 25584 37179 25642 37185
rect 25584 37145 25596 37179
rect 25630 37176 25642 37179
rect 26602 37176 26608 37188
rect 25630 37148 26608 37176
rect 25630 37145 25642 37148
rect 25584 37139 25642 37145
rect 26602 37136 26608 37148
rect 26660 37136 26666 37188
rect 22922 37108 22928 37120
rect 22020 37080 22928 37108
rect 22922 37068 22928 37080
rect 22980 37068 22986 37120
rect 24854 37108 24860 37120
rect 24815 37080 24860 37108
rect 24854 37068 24860 37080
rect 24912 37068 24918 37120
rect 25498 37068 25504 37120
rect 25556 37068 25562 37120
rect 27356 37108 27384 37207
rect 28074 37204 28080 37256
rect 28132 37244 28138 37256
rect 28350 37244 28356 37256
rect 28132 37216 28177 37244
rect 28311 37216 28356 37244
rect 28132 37204 28138 37216
rect 28350 37204 28356 37216
rect 28408 37204 28414 37256
rect 30006 37244 30012 37256
rect 29967 37216 30012 37244
rect 30006 37204 30012 37216
rect 30064 37204 30070 37256
rect 32766 37244 32772 37256
rect 32727 37216 32772 37244
rect 32766 37204 32772 37216
rect 32824 37204 32830 37256
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 33560 37216 34897 37244
rect 33560 37204 33566 37216
rect 34885 37213 34897 37216
rect 34931 37213 34943 37247
rect 34885 37207 34943 37213
rect 35713 37247 35771 37253
rect 35713 37213 35725 37247
rect 35759 37244 35771 37247
rect 35802 37244 35808 37256
rect 35759 37216 35808 37244
rect 35759 37213 35771 37216
rect 35713 37207 35771 37213
rect 35802 37204 35808 37216
rect 35860 37204 35866 37256
rect 36740 37253 36768 37284
rect 39114 37272 39120 37284
rect 39172 37312 39178 37324
rect 39172 37284 39528 37312
rect 39172 37272 39178 37284
rect 39500 37256 39528 37284
rect 39574 37272 39580 37324
rect 39632 37312 39638 37324
rect 41141 37315 41199 37321
rect 39632 37284 41092 37312
rect 39632 37272 39638 37284
rect 36725 37247 36783 37253
rect 36725 37213 36737 37247
rect 36771 37213 36783 37247
rect 38930 37244 38936 37256
rect 38891 37216 38936 37244
rect 36725 37207 36783 37213
rect 38930 37204 38936 37216
rect 38988 37204 38994 37256
rect 39022 37204 39028 37256
rect 39080 37244 39086 37256
rect 39209 37247 39267 37253
rect 39080 37216 39125 37244
rect 39080 37204 39086 37216
rect 39209 37213 39221 37247
rect 39255 37244 39267 37247
rect 39390 37244 39396 37256
rect 39255 37216 39396 37244
rect 39255 37213 39267 37216
rect 39209 37207 39267 37213
rect 39390 37204 39396 37216
rect 39448 37204 39454 37256
rect 39482 37204 39488 37256
rect 39540 37204 39546 37256
rect 40862 37204 40868 37256
rect 40920 37244 40926 37256
rect 40957 37247 41015 37253
rect 40957 37244 40969 37247
rect 40920 37216 40969 37244
rect 40920 37204 40926 37216
rect 40957 37213 40969 37216
rect 41003 37213 41015 37247
rect 41064 37244 41092 37284
rect 41141 37281 41153 37315
rect 41187 37312 41199 37315
rect 41386 37312 41414 37352
rect 43070 37340 43076 37352
rect 43128 37340 43134 37392
rect 41601 37315 41659 37321
rect 41601 37312 41613 37315
rect 41187 37284 41414 37312
rect 41524 37284 41613 37312
rect 41187 37281 41199 37284
rect 41141 37275 41199 37281
rect 41524 37244 41552 37284
rect 41601 37281 41613 37284
rect 41647 37312 41659 37315
rect 41647 37284 43024 37312
rect 41647 37281 41659 37284
rect 41601 37275 41659 37281
rect 41874 37244 41880 37256
rect 41064 37216 41552 37244
rect 41835 37216 41880 37244
rect 40957 37207 41015 37213
rect 41874 37204 41880 37216
rect 41932 37244 41938 37256
rect 42794 37244 42800 37256
rect 41932 37216 42800 37244
rect 41932 37204 41938 37216
rect 42794 37204 42800 37216
rect 42852 37204 42858 37256
rect 42996 37253 43024 37284
rect 42981 37247 43039 37253
rect 42981 37213 42993 37247
rect 43027 37213 43039 37247
rect 42981 37207 43039 37213
rect 44085 37247 44143 37253
rect 44085 37213 44097 37247
rect 44131 37244 44143 37247
rect 44358 37244 44364 37256
rect 44131 37216 44364 37244
rect 44131 37213 44143 37216
rect 44085 37207 44143 37213
rect 44358 37204 44364 37216
rect 44416 37204 44422 37256
rect 45186 37244 45192 37256
rect 45147 37216 45192 37244
rect 45186 37204 45192 37216
rect 45244 37204 45250 37256
rect 46842 37204 46848 37256
rect 46900 37244 46906 37256
rect 47213 37247 47271 37253
rect 47213 37244 47225 37247
rect 46900 37216 47225 37244
rect 46900 37204 46906 37216
rect 47213 37213 47225 37216
rect 47259 37213 47271 37247
rect 47213 37207 47271 37213
rect 33036 37179 33094 37185
rect 33036 37145 33048 37179
rect 33082 37176 33094 37179
rect 43165 37179 43223 37185
rect 33082 37148 34744 37176
rect 33082 37145 33094 37148
rect 33036 37139 33094 37145
rect 29822 37108 29828 37120
rect 27356 37080 29828 37108
rect 29822 37068 29828 37080
rect 29880 37108 29886 37120
rect 30374 37108 30380 37120
rect 29880 37080 30380 37108
rect 29880 37068 29886 37080
rect 30374 37068 30380 37080
rect 30432 37068 30438 37120
rect 33870 37068 33876 37120
rect 33928 37108 33934 37120
rect 34716 37117 34744 37148
rect 43165 37145 43177 37179
rect 43211 37176 43223 37179
rect 43254 37176 43260 37188
rect 43211 37148 43260 37176
rect 43211 37145 43223 37148
rect 43165 37139 43223 37145
rect 43254 37136 43260 37148
rect 43312 37136 43318 37188
rect 44269 37179 44327 37185
rect 44269 37145 44281 37179
rect 44315 37176 44327 37179
rect 44726 37176 44732 37188
rect 44315 37148 44732 37176
rect 44315 37145 44327 37148
rect 44269 37139 44327 37145
rect 44726 37136 44732 37148
rect 44784 37136 44790 37188
rect 44818 37136 44824 37188
rect 44876 37176 44882 37188
rect 45434 37179 45492 37185
rect 45434 37176 45446 37179
rect 44876 37148 45446 37176
rect 44876 37136 44882 37148
rect 45434 37145 45446 37148
rect 45480 37145 45492 37179
rect 45434 37139 45492 37145
rect 34149 37111 34207 37117
rect 34149 37108 34161 37111
rect 33928 37080 34161 37108
rect 33928 37068 33934 37080
rect 34149 37077 34161 37080
rect 34195 37077 34207 37111
rect 34149 37071 34207 37077
rect 34701 37111 34759 37117
rect 34701 37077 34713 37111
rect 34747 37077 34759 37111
rect 34701 37071 34759 37077
rect 35986 37068 35992 37120
rect 36044 37108 36050 37120
rect 36909 37111 36967 37117
rect 36909 37108 36921 37111
rect 36044 37080 36921 37108
rect 36044 37068 36050 37080
rect 36909 37077 36921 37080
rect 36955 37077 36967 37111
rect 36909 37071 36967 37077
rect 45002 37068 45008 37120
rect 45060 37108 45066 37120
rect 46566 37108 46572 37120
rect 45060 37080 46572 37108
rect 45060 37068 45066 37080
rect 46566 37068 46572 37080
rect 46624 37068 46630 37120
rect 1104 37018 68816 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 68816 37018
rect 1104 36944 68816 36966
rect 22738 36904 22744 36916
rect 22699 36876 22744 36904
rect 22738 36864 22744 36876
rect 22796 36864 22802 36916
rect 24670 36904 24676 36916
rect 24631 36876 24676 36904
rect 24670 36864 24676 36876
rect 24728 36864 24734 36916
rect 29730 36864 29736 36916
rect 29788 36904 29794 36916
rect 30006 36904 30012 36916
rect 30064 36913 30070 36916
rect 30064 36907 30083 36913
rect 29788 36876 30012 36904
rect 29788 36864 29794 36876
rect 30006 36864 30012 36876
rect 30071 36873 30083 36907
rect 30190 36904 30196 36916
rect 30151 36876 30196 36904
rect 30064 36867 30083 36873
rect 30064 36864 30070 36867
rect 30190 36864 30196 36876
rect 30248 36864 30254 36916
rect 37826 36904 37832 36916
rect 34072 36876 36216 36904
rect 25682 36836 25688 36848
rect 6886 36808 25688 36836
rect 2501 36771 2559 36777
rect 2501 36737 2513 36771
rect 2547 36768 2559 36771
rect 6886 36768 6914 36808
rect 25682 36796 25688 36808
rect 25740 36796 25746 36848
rect 29822 36836 29828 36848
rect 29783 36808 29828 36836
rect 29822 36796 29828 36808
rect 29880 36796 29886 36848
rect 32674 36836 32680 36848
rect 29932 36808 32680 36836
rect 2547 36740 6914 36768
rect 22649 36771 22707 36777
rect 2547 36737 2559 36740
rect 2501 36731 2559 36737
rect 22649 36737 22661 36771
rect 22695 36737 22707 36771
rect 22649 36731 22707 36737
rect 22664 36700 22692 36731
rect 23290 36728 23296 36780
rect 23348 36768 23354 36780
rect 23385 36771 23443 36777
rect 23385 36768 23397 36771
rect 23348 36740 23397 36768
rect 23348 36728 23354 36740
rect 23385 36737 23397 36740
rect 23431 36737 23443 36771
rect 24854 36768 24860 36780
rect 24815 36740 24860 36768
rect 23385 36731 23443 36737
rect 24854 36728 24860 36740
rect 24912 36728 24918 36780
rect 25498 36728 25504 36780
rect 25556 36768 25562 36780
rect 25869 36771 25927 36777
rect 25869 36768 25881 36771
rect 25556 36740 25881 36768
rect 25556 36728 25562 36740
rect 25869 36737 25881 36740
rect 25915 36737 25927 36771
rect 25869 36731 25927 36737
rect 27249 36771 27307 36777
rect 27249 36737 27261 36771
rect 27295 36768 27307 36771
rect 27295 36766 29792 36768
rect 29932 36766 29960 36808
rect 32674 36796 32680 36808
rect 32732 36796 32738 36848
rect 27295 36740 29960 36766
rect 27295 36737 27307 36740
rect 29764 36738 29960 36740
rect 27249 36731 27307 36737
rect 30190 36728 30196 36780
rect 30248 36768 30254 36780
rect 30745 36771 30803 36777
rect 30745 36768 30757 36771
rect 30248 36740 30757 36768
rect 30248 36728 30254 36740
rect 30745 36737 30757 36740
rect 30791 36737 30803 36771
rect 32585 36771 32643 36777
rect 32585 36768 32597 36771
rect 30745 36731 30803 36737
rect 31726 36740 32597 36768
rect 25593 36703 25651 36709
rect 22664 36672 23704 36700
rect 1578 36524 1584 36576
rect 1636 36564 1642 36576
rect 23676 36573 23704 36672
rect 25593 36669 25605 36703
rect 25639 36700 25651 36703
rect 26234 36700 26240 36712
rect 25639 36672 26240 36700
rect 25639 36669 25651 36672
rect 25593 36663 25651 36669
rect 26234 36660 26240 36672
rect 26292 36700 26298 36712
rect 26292 36672 27292 36700
rect 26292 36660 26298 36672
rect 2593 36567 2651 36573
rect 2593 36564 2605 36567
rect 1636 36536 2605 36564
rect 1636 36524 1642 36536
rect 2593 36533 2605 36536
rect 2639 36533 2651 36567
rect 2593 36527 2651 36533
rect 23661 36567 23719 36573
rect 23661 36533 23673 36567
rect 23707 36564 23719 36567
rect 24302 36564 24308 36576
rect 23707 36536 24308 36564
rect 23707 36533 23719 36536
rect 23661 36527 23719 36533
rect 24302 36524 24308 36536
rect 24360 36524 24366 36576
rect 27264 36564 27292 36672
rect 27338 36660 27344 36712
rect 27396 36700 27402 36712
rect 27525 36703 27583 36709
rect 27525 36700 27537 36703
rect 27396 36672 27537 36700
rect 27396 36660 27402 36672
rect 27525 36669 27537 36672
rect 27571 36669 27583 36703
rect 27525 36663 27583 36669
rect 28537 36703 28595 36709
rect 28537 36669 28549 36703
rect 28583 36669 28595 36703
rect 28810 36700 28816 36712
rect 28771 36672 28816 36700
rect 28537 36663 28595 36669
rect 28552 36632 28580 36663
rect 28810 36660 28816 36672
rect 28868 36660 28874 36712
rect 31021 36703 31079 36709
rect 31021 36669 31033 36703
rect 31067 36700 31079 36703
rect 31386 36700 31392 36712
rect 31067 36672 31392 36700
rect 31067 36669 31079 36672
rect 31021 36663 31079 36669
rect 31386 36660 31392 36672
rect 31444 36660 31450 36712
rect 29546 36632 29552 36644
rect 28552 36604 29552 36632
rect 29546 36592 29552 36604
rect 29604 36632 29610 36644
rect 31726 36632 31754 36740
rect 32585 36737 32597 36740
rect 32631 36737 32643 36771
rect 32585 36731 32643 36737
rect 32861 36771 32919 36777
rect 32861 36737 32873 36771
rect 32907 36768 32919 36771
rect 33318 36768 33324 36780
rect 32907 36740 33324 36768
rect 32907 36737 32919 36740
rect 32861 36731 32919 36737
rect 33318 36728 33324 36740
rect 33376 36728 33382 36780
rect 33870 36768 33876 36780
rect 33831 36740 33876 36768
rect 33870 36728 33876 36740
rect 33928 36728 33934 36780
rect 34072 36777 34100 36876
rect 36188 36848 36216 36876
rect 37568 36876 37832 36904
rect 36170 36836 36176 36848
rect 36083 36808 36176 36836
rect 36170 36796 36176 36808
rect 36228 36796 36234 36848
rect 37568 36845 37596 36876
rect 37826 36864 37832 36876
rect 37884 36904 37890 36916
rect 38378 36904 38384 36916
rect 37884 36876 38384 36904
rect 37884 36864 37890 36876
rect 38378 36864 38384 36876
rect 38436 36864 38442 36916
rect 38930 36864 38936 36916
rect 38988 36904 38994 36916
rect 39393 36907 39451 36913
rect 39393 36904 39405 36907
rect 38988 36876 39405 36904
rect 38988 36864 38994 36876
rect 39393 36873 39405 36876
rect 39439 36873 39451 36907
rect 39393 36867 39451 36873
rect 39592 36876 42288 36904
rect 36373 36839 36431 36845
rect 36373 36836 36385 36839
rect 36280 36808 36385 36836
rect 34057 36771 34115 36777
rect 34057 36737 34069 36771
rect 34103 36737 34115 36771
rect 34057 36731 34115 36737
rect 35802 36728 35808 36780
rect 35860 36768 35866 36780
rect 36280 36768 36308 36808
rect 36373 36805 36385 36808
rect 36419 36805 36431 36839
rect 36373 36799 36431 36805
rect 37553 36839 37611 36845
rect 37553 36805 37565 36839
rect 37599 36805 37611 36839
rect 37553 36799 37611 36805
rect 37737 36839 37795 36845
rect 37737 36805 37749 36839
rect 37783 36836 37795 36839
rect 39592 36836 39620 36876
rect 37783 36808 39620 36836
rect 37783 36805 37795 36808
rect 37737 36799 37795 36805
rect 40586 36796 40592 36848
rect 40644 36836 40650 36848
rect 40681 36839 40739 36845
rect 40681 36836 40693 36839
rect 40644 36808 40693 36836
rect 40644 36796 40650 36808
rect 40681 36805 40693 36808
rect 40727 36805 40739 36839
rect 40681 36799 40739 36805
rect 37366 36768 37372 36780
rect 35860 36740 36308 36768
rect 37327 36740 37372 36768
rect 35860 36728 35866 36740
rect 37366 36728 37372 36740
rect 37424 36728 37430 36780
rect 38197 36771 38255 36777
rect 38197 36737 38209 36771
rect 38243 36737 38255 36771
rect 38378 36768 38384 36780
rect 38339 36740 38384 36768
rect 38197 36731 38255 36737
rect 34790 36700 34796 36712
rect 34751 36672 34796 36700
rect 34790 36660 34796 36672
rect 34848 36660 34854 36712
rect 34882 36660 34888 36712
rect 34940 36709 34946 36712
rect 34940 36703 34968 36709
rect 34956 36669 34968 36703
rect 34940 36663 34968 36669
rect 35069 36703 35127 36709
rect 35069 36669 35081 36703
rect 35115 36700 35127 36703
rect 35434 36700 35440 36712
rect 35115 36672 35440 36700
rect 35115 36669 35127 36672
rect 35069 36663 35127 36669
rect 34940 36660 34946 36663
rect 35434 36660 35440 36672
rect 35492 36660 35498 36712
rect 35713 36703 35771 36709
rect 35713 36669 35725 36703
rect 35759 36700 35771 36703
rect 38212 36700 38240 36731
rect 38378 36728 38384 36740
rect 38436 36728 38442 36780
rect 39022 36768 39028 36780
rect 38983 36740 39028 36768
rect 39022 36728 39028 36740
rect 39080 36728 39086 36780
rect 39206 36768 39212 36780
rect 39167 36740 39212 36768
rect 39206 36728 39212 36740
rect 39264 36728 39270 36780
rect 41601 36771 41659 36777
rect 41601 36768 41613 36771
rect 41386 36740 41613 36768
rect 35759 36672 38240 36700
rect 38565 36703 38623 36709
rect 35759 36669 35771 36672
rect 35713 36663 35771 36669
rect 38565 36669 38577 36703
rect 38611 36700 38623 36703
rect 41386 36700 41414 36740
rect 41601 36737 41613 36740
rect 41647 36737 41659 36771
rect 41601 36731 41659 36737
rect 41693 36771 41751 36777
rect 41693 36737 41705 36771
rect 41739 36768 41751 36771
rect 41874 36768 41880 36780
rect 41739 36740 41880 36768
rect 41739 36737 41751 36740
rect 41693 36731 41751 36737
rect 41874 36728 41880 36740
rect 41932 36728 41938 36780
rect 42260 36768 42288 36876
rect 42702 36864 42708 36916
rect 42760 36904 42766 36916
rect 43346 36904 43352 36916
rect 42760 36876 43352 36904
rect 42760 36864 42766 36876
rect 43346 36864 43352 36876
rect 43404 36864 43410 36916
rect 44818 36904 44824 36916
rect 44779 36876 44824 36904
rect 44818 36864 44824 36876
rect 44876 36864 44882 36916
rect 44910 36864 44916 36916
rect 44968 36904 44974 36916
rect 45370 36904 45376 36916
rect 44968 36876 45376 36904
rect 44968 36864 44974 36876
rect 45370 36864 45376 36876
rect 45428 36904 45434 36916
rect 45428 36876 46336 36904
rect 45428 36864 45434 36876
rect 42426 36796 42432 36848
rect 42484 36836 42490 36848
rect 43901 36839 43959 36845
rect 43901 36836 43913 36839
rect 42484 36808 43913 36836
rect 42484 36796 42490 36808
rect 43901 36805 43913 36808
rect 43947 36805 43959 36839
rect 43901 36799 43959 36805
rect 43165 36771 43223 36777
rect 43165 36768 43177 36771
rect 42260 36740 43177 36768
rect 43165 36737 43177 36740
rect 43211 36737 43223 36771
rect 43165 36731 43223 36737
rect 43254 36728 43260 36780
rect 43312 36768 43318 36780
rect 44085 36771 44143 36777
rect 43312 36740 43357 36768
rect 43312 36728 43318 36740
rect 44085 36737 44097 36771
rect 44131 36768 44143 36771
rect 44818 36768 44824 36780
rect 44131 36740 44824 36768
rect 44131 36737 44143 36740
rect 44085 36731 44143 36737
rect 44818 36728 44824 36740
rect 44876 36728 44882 36780
rect 45077 36771 45135 36777
rect 45077 36737 45089 36771
rect 45123 36768 45135 36771
rect 45170 36774 45228 36780
rect 45123 36737 45140 36768
rect 45077 36731 45140 36737
rect 45170 36740 45182 36774
rect 45216 36771 45228 36774
rect 45270 36771 45328 36777
rect 45216 36768 45229 36771
rect 45216 36740 45232 36768
rect 45170 36734 45232 36740
rect 38611 36672 41414 36700
rect 41509 36703 41567 36709
rect 38611 36669 38623 36672
rect 38565 36663 38623 36669
rect 41509 36669 41521 36703
rect 41555 36669 41567 36703
rect 41509 36663 41567 36669
rect 41785 36703 41843 36709
rect 41785 36669 41797 36703
rect 41831 36700 41843 36703
rect 42702 36700 42708 36712
rect 41831 36672 42708 36700
rect 41831 36669 41843 36672
rect 41785 36663 41843 36669
rect 34514 36632 34520 36644
rect 29604 36604 31754 36632
rect 34475 36604 34520 36632
rect 29604 36592 29610 36604
rect 34514 36592 34520 36604
rect 34572 36592 34578 36644
rect 41524 36632 41552 36663
rect 42702 36660 42708 36672
rect 42760 36660 42766 36712
rect 43073 36703 43131 36709
rect 43073 36669 43085 36703
rect 43119 36700 43131 36703
rect 43346 36700 43352 36712
rect 43119 36672 43208 36700
rect 43307 36672 43352 36700
rect 43119 36669 43131 36672
rect 43073 36663 43131 36669
rect 42794 36632 42800 36644
rect 41524 36604 42800 36632
rect 42794 36592 42800 36604
rect 42852 36592 42858 36644
rect 43180 36632 43208 36672
rect 43346 36660 43352 36672
rect 43404 36660 43410 36712
rect 44910 36660 44916 36712
rect 44968 36700 44974 36712
rect 45112 36700 45140 36731
rect 44968 36672 45140 36700
rect 44968 36660 44974 36672
rect 45204 36644 45232 36734
rect 45270 36737 45282 36771
rect 45316 36737 45328 36771
rect 45270 36731 45328 36737
rect 45465 36771 45523 36777
rect 45465 36737 45477 36771
rect 45511 36768 45523 36771
rect 45646 36768 45652 36780
rect 45511 36740 45652 36768
rect 45511 36737 45523 36740
rect 45465 36731 45523 36737
rect 44269 36635 44327 36641
rect 44269 36632 44281 36635
rect 43180 36604 44281 36632
rect 44269 36601 44281 36604
rect 44315 36601 44327 36635
rect 44269 36595 44327 36601
rect 44726 36592 44732 36644
rect 44784 36632 44790 36644
rect 45186 36632 45192 36644
rect 44784 36604 45192 36632
rect 44784 36592 44790 36604
rect 45186 36592 45192 36604
rect 45244 36592 45250 36644
rect 29914 36564 29920 36576
rect 27264 36536 29920 36564
rect 29914 36524 29920 36536
rect 29972 36524 29978 36576
rect 30009 36567 30067 36573
rect 30009 36533 30021 36567
rect 30055 36564 30067 36567
rect 30466 36564 30472 36576
rect 30055 36536 30472 36564
rect 30055 36533 30067 36536
rect 30009 36527 30067 36533
rect 30466 36524 30472 36536
rect 30524 36524 30530 36576
rect 35526 36524 35532 36576
rect 35584 36564 35590 36576
rect 35710 36564 35716 36576
rect 35584 36536 35716 36564
rect 35584 36524 35590 36536
rect 35710 36524 35716 36536
rect 35768 36564 35774 36576
rect 36357 36567 36415 36573
rect 36357 36564 36369 36567
rect 35768 36536 36369 36564
rect 35768 36524 35774 36536
rect 36357 36533 36369 36536
rect 36403 36533 36415 36567
rect 36538 36564 36544 36576
rect 36499 36536 36544 36564
rect 36357 36527 36415 36533
rect 36538 36524 36544 36536
rect 36596 36524 36602 36576
rect 40402 36524 40408 36576
rect 40460 36564 40466 36576
rect 40773 36567 40831 36573
rect 40773 36564 40785 36567
rect 40460 36536 40785 36564
rect 40460 36524 40466 36536
rect 40773 36533 40785 36536
rect 40819 36533 40831 36567
rect 41322 36564 41328 36576
rect 41283 36536 41328 36564
rect 40773 36527 40831 36533
rect 41322 36524 41328 36536
rect 41380 36524 41386 36576
rect 42889 36567 42947 36573
rect 42889 36533 42901 36567
rect 42935 36564 42947 36567
rect 45296 36564 45324 36731
rect 45646 36728 45652 36740
rect 45704 36768 45710 36780
rect 46308 36777 46336 36876
rect 46201 36771 46259 36777
rect 45704 36740 45968 36768
rect 45704 36728 45710 36740
rect 45940 36632 45968 36740
rect 46201 36737 46213 36771
rect 46247 36737 46259 36771
rect 46201 36731 46259 36737
rect 46293 36771 46351 36777
rect 46293 36737 46305 36771
rect 46339 36737 46351 36771
rect 46293 36731 46351 36737
rect 46216 36700 46244 36731
rect 46382 36728 46388 36780
rect 46440 36768 46446 36780
rect 46569 36771 46627 36777
rect 46440 36740 46485 36768
rect 46440 36728 46446 36740
rect 46569 36737 46581 36771
rect 46615 36768 46627 36771
rect 46750 36768 46756 36780
rect 46615 36740 46756 36768
rect 46615 36737 46627 36740
rect 46569 36731 46627 36737
rect 46750 36728 46756 36740
rect 46808 36728 46814 36780
rect 47854 36700 47860 36712
rect 46216 36672 47860 36700
rect 47854 36660 47860 36672
rect 47912 36660 47918 36712
rect 46750 36632 46756 36644
rect 45940 36604 46756 36632
rect 46750 36592 46756 36604
rect 46808 36592 46814 36644
rect 42935 36536 45324 36564
rect 45925 36567 45983 36573
rect 42935 36533 42947 36536
rect 42889 36527 42947 36533
rect 45925 36533 45937 36567
rect 45971 36564 45983 36567
rect 46566 36564 46572 36576
rect 45971 36536 46572 36564
rect 45971 36533 45983 36536
rect 45925 36527 45983 36533
rect 46566 36524 46572 36536
rect 46624 36524 46630 36576
rect 1104 36474 68816 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 68816 36474
rect 1104 36400 68816 36422
rect 26602 36360 26608 36372
rect 26563 36332 26608 36360
rect 26602 36320 26608 36332
rect 26660 36320 26666 36372
rect 32306 36360 32312 36372
rect 32267 36332 32312 36360
rect 32306 36320 32312 36332
rect 32364 36320 32370 36372
rect 33226 36320 33232 36372
rect 33284 36360 33290 36372
rect 33321 36363 33379 36369
rect 33321 36360 33333 36363
rect 33284 36332 33333 36360
rect 33284 36320 33290 36332
rect 33321 36329 33333 36332
rect 33367 36329 33379 36363
rect 33502 36360 33508 36372
rect 33463 36332 33508 36360
rect 33321 36323 33379 36329
rect 33502 36320 33508 36332
rect 33560 36320 33566 36372
rect 36170 36320 36176 36372
rect 36228 36360 36234 36372
rect 37369 36363 37427 36369
rect 37369 36360 37381 36363
rect 36228 36332 37381 36360
rect 36228 36320 36234 36332
rect 37369 36329 37381 36332
rect 37415 36329 37427 36363
rect 37369 36323 37427 36329
rect 39206 36320 39212 36372
rect 39264 36360 39270 36372
rect 39301 36363 39359 36369
rect 39301 36360 39313 36363
rect 39264 36332 39313 36360
rect 39264 36320 39270 36332
rect 39301 36329 39313 36332
rect 39347 36329 39359 36363
rect 39301 36323 39359 36329
rect 41322 36320 41328 36372
rect 41380 36360 41386 36372
rect 46382 36360 46388 36372
rect 41380 36332 46388 36360
rect 41380 36320 41386 36332
rect 46382 36320 46388 36332
rect 46440 36320 46446 36372
rect 47854 36360 47860 36372
rect 47815 36332 47860 36360
rect 47854 36320 47860 36332
rect 47912 36320 47918 36372
rect 23661 36295 23719 36301
rect 23661 36261 23673 36295
rect 23707 36261 23719 36295
rect 23661 36255 23719 36261
rect 1578 36224 1584 36236
rect 1539 36196 1584 36224
rect 1578 36184 1584 36196
rect 1636 36184 1642 36236
rect 2774 36224 2780 36236
rect 2735 36196 2780 36224
rect 2774 36184 2780 36196
rect 2832 36184 2838 36236
rect 23676 36224 23704 36255
rect 24397 36227 24455 36233
rect 24397 36224 24409 36227
rect 23676 36196 24409 36224
rect 24397 36193 24409 36196
rect 24443 36224 24455 36227
rect 28074 36224 28080 36236
rect 24443 36196 28080 36224
rect 24443 36193 24455 36196
rect 24397 36187 24455 36193
rect 28074 36184 28080 36196
rect 28132 36184 28138 36236
rect 30834 36224 30840 36236
rect 30300 36196 30840 36224
rect 1394 36156 1400 36168
rect 1355 36128 1400 36156
rect 1394 36116 1400 36128
rect 1452 36116 1458 36168
rect 22278 36156 22284 36168
rect 22239 36128 22284 36156
rect 22278 36116 22284 36128
rect 22336 36116 22342 36168
rect 23566 36116 23572 36168
rect 23624 36156 23630 36168
rect 24581 36159 24639 36165
rect 24581 36156 24593 36159
rect 23624 36128 24593 36156
rect 23624 36116 23630 36128
rect 24581 36125 24593 36128
rect 24627 36125 24639 36159
rect 24581 36119 24639 36125
rect 25225 36159 25283 36165
rect 25225 36125 25237 36159
rect 25271 36156 25283 36159
rect 25774 36156 25780 36168
rect 25271 36128 25780 36156
rect 25271 36125 25283 36128
rect 25225 36119 25283 36125
rect 25774 36116 25780 36128
rect 25832 36116 25838 36168
rect 26789 36159 26847 36165
rect 26789 36125 26801 36159
rect 26835 36156 26847 36159
rect 27522 36156 27528 36168
rect 26835 36128 27528 36156
rect 26835 36125 26847 36128
rect 26789 36119 26847 36125
rect 27522 36116 27528 36128
rect 27580 36116 27586 36168
rect 28442 36116 28448 36168
rect 28500 36156 28506 36168
rect 28537 36159 28595 36165
rect 28537 36156 28549 36159
rect 28500 36128 28549 36156
rect 28500 36116 28506 36128
rect 28537 36125 28549 36128
rect 28583 36125 28595 36159
rect 28537 36119 28595 36125
rect 29733 36159 29791 36165
rect 29733 36125 29745 36159
rect 29779 36156 29791 36159
rect 29914 36156 29920 36168
rect 29779 36128 29920 36156
rect 29779 36125 29791 36128
rect 29733 36119 29791 36125
rect 22548 36091 22606 36097
rect 22548 36057 22560 36091
rect 22594 36088 22606 36091
rect 23014 36088 23020 36100
rect 22594 36060 23020 36088
rect 22594 36057 22606 36060
rect 22548 36051 22606 36057
rect 23014 36048 23020 36060
rect 23072 36048 23078 36100
rect 28552 36088 28580 36119
rect 29914 36116 29920 36128
rect 29972 36116 29978 36168
rect 30300 36165 30328 36196
rect 30834 36184 30840 36196
rect 30892 36184 30898 36236
rect 35986 36224 35992 36236
rect 35947 36196 35992 36224
rect 35986 36184 35992 36196
rect 36044 36184 36050 36236
rect 39022 36184 39028 36236
rect 39080 36224 39086 36236
rect 40129 36227 40187 36233
rect 40129 36224 40141 36227
rect 39080 36196 40141 36224
rect 39080 36184 39086 36196
rect 40129 36193 40141 36196
rect 40175 36193 40187 36227
rect 40129 36187 40187 36193
rect 43349 36227 43407 36233
rect 43349 36193 43361 36227
rect 43395 36224 43407 36227
rect 44818 36224 44824 36236
rect 43395 36196 44824 36224
rect 43395 36193 43407 36196
rect 43349 36187 43407 36193
rect 44818 36184 44824 36196
rect 44876 36184 44882 36236
rect 30285 36159 30343 36165
rect 30285 36125 30297 36159
rect 30331 36125 30343 36159
rect 30285 36119 30343 36125
rect 30469 36159 30527 36165
rect 30469 36125 30481 36159
rect 30515 36156 30527 36159
rect 30929 36159 30987 36165
rect 30929 36156 30941 36159
rect 30515 36128 30941 36156
rect 30515 36125 30527 36128
rect 30469 36119 30527 36125
rect 30929 36125 30941 36128
rect 30975 36125 30987 36159
rect 34698 36156 34704 36168
rect 30929 36119 30987 36125
rect 31036 36128 34704 36156
rect 31036 36088 31064 36128
rect 34698 36116 34704 36128
rect 34756 36116 34762 36168
rect 37918 36156 37924 36168
rect 37879 36128 37924 36156
rect 37918 36116 37924 36128
rect 37976 36116 37982 36168
rect 39758 36116 39764 36168
rect 39816 36156 39822 36168
rect 39853 36159 39911 36165
rect 39853 36156 39865 36159
rect 39816 36128 39865 36156
rect 39816 36116 39822 36128
rect 39853 36125 39865 36128
rect 39899 36156 39911 36159
rect 41509 36159 41567 36165
rect 41509 36156 41521 36159
rect 39899 36128 41521 36156
rect 39899 36125 39911 36128
rect 39853 36119 39911 36125
rect 41509 36125 41521 36128
rect 41555 36125 41567 36159
rect 41509 36119 41567 36125
rect 41785 36159 41843 36165
rect 41785 36125 41797 36159
rect 41831 36156 41843 36159
rect 42426 36156 42432 36168
rect 41831 36128 42432 36156
rect 41831 36125 41843 36128
rect 41785 36119 41843 36125
rect 42426 36116 42432 36128
rect 42484 36116 42490 36168
rect 42978 36116 42984 36168
rect 43036 36156 43042 36168
rect 43533 36159 43591 36165
rect 43533 36156 43545 36159
rect 43036 36128 43545 36156
rect 43036 36116 43042 36128
rect 43533 36125 43545 36128
rect 43579 36125 43591 36159
rect 43533 36119 43591 36125
rect 45554 36116 45560 36168
rect 45612 36156 45618 36168
rect 46477 36159 46535 36165
rect 46477 36156 46489 36159
rect 45612 36128 46489 36156
rect 45612 36116 45618 36128
rect 46477 36125 46489 36128
rect 46523 36125 46535 36159
rect 46477 36119 46535 36125
rect 46566 36116 46572 36168
rect 46624 36156 46630 36168
rect 46733 36159 46791 36165
rect 46733 36156 46745 36159
rect 46624 36128 46745 36156
rect 46624 36116 46630 36128
rect 46733 36125 46745 36128
rect 46779 36125 46791 36159
rect 46733 36119 46791 36125
rect 66898 36116 66904 36168
rect 66956 36156 66962 36168
rect 67913 36159 67971 36165
rect 67913 36156 67925 36159
rect 66956 36128 67925 36156
rect 66956 36116 66962 36128
rect 67913 36125 67925 36128
rect 67959 36125 67971 36159
rect 67913 36119 67971 36125
rect 28552 36060 31064 36088
rect 31196 36091 31254 36097
rect 31196 36057 31208 36091
rect 31242 36088 31254 36091
rect 31294 36088 31300 36100
rect 31242 36060 31300 36088
rect 31242 36057 31254 36060
rect 31196 36051 31254 36057
rect 31294 36048 31300 36060
rect 31352 36048 31358 36100
rect 33137 36091 33195 36097
rect 33137 36057 33149 36091
rect 33183 36088 33195 36091
rect 33870 36088 33876 36100
rect 33183 36060 33876 36088
rect 33183 36057 33195 36060
rect 33137 36051 33195 36057
rect 33870 36048 33876 36060
rect 33928 36048 33934 36100
rect 36256 36091 36314 36097
rect 36256 36057 36268 36091
rect 36302 36088 36314 36091
rect 36354 36088 36360 36100
rect 36302 36060 36360 36088
rect 36302 36057 36314 36060
rect 36256 36051 36314 36057
rect 36354 36048 36360 36060
rect 36412 36048 36418 36100
rect 38188 36091 38246 36097
rect 38188 36057 38200 36091
rect 38234 36088 38246 36091
rect 38930 36088 38936 36100
rect 38234 36060 38936 36088
rect 38234 36057 38246 36060
rect 38188 36051 38246 36057
rect 38930 36048 38936 36060
rect 38988 36048 38994 36100
rect 23750 35980 23756 36032
rect 23808 36020 23814 36032
rect 24765 36023 24823 36029
rect 24765 36020 24777 36023
rect 23808 35992 24777 36020
rect 23808 35980 23814 35992
rect 24765 35989 24777 35992
rect 24811 35989 24823 36023
rect 25314 36020 25320 36032
rect 25275 35992 25320 36020
rect 24765 35983 24823 35989
rect 25314 35980 25320 35992
rect 25372 35980 25378 36032
rect 28718 36020 28724 36032
rect 28679 35992 28724 36020
rect 28718 35980 28724 35992
rect 28776 35980 28782 36032
rect 29546 36020 29552 36032
rect 29507 35992 29552 36020
rect 29546 35980 29552 35992
rect 29604 35980 29610 36032
rect 33318 35980 33324 36032
rect 33376 36029 33382 36032
rect 33376 36023 33395 36029
rect 33383 35989 33395 36023
rect 33376 35983 33395 35989
rect 43717 36023 43775 36029
rect 43717 35989 43729 36023
rect 43763 36020 43775 36023
rect 44174 36020 44180 36032
rect 43763 35992 44180 36020
rect 43763 35989 43775 35992
rect 43717 35983 43775 35989
rect 33376 35980 33382 35983
rect 44174 35980 44180 35992
rect 44232 35980 44238 36032
rect 1104 35930 68816 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 68816 35930
rect 1104 35856 68816 35878
rect 19705 35819 19763 35825
rect 19705 35785 19717 35819
rect 19751 35816 19763 35819
rect 23201 35819 23259 35825
rect 19751 35788 23060 35816
rect 19751 35785 19763 35788
rect 19705 35779 19763 35785
rect 14458 35708 14464 35760
rect 14516 35748 14522 35760
rect 20073 35751 20131 35757
rect 20073 35748 20085 35751
rect 14516 35720 20085 35748
rect 14516 35708 14522 35720
rect 20073 35717 20085 35720
rect 20119 35748 20131 35751
rect 20119 35720 21036 35748
rect 20119 35717 20131 35720
rect 20073 35711 20131 35717
rect 1394 35640 1400 35692
rect 1452 35680 1458 35692
rect 2133 35683 2191 35689
rect 2133 35680 2145 35683
rect 1452 35652 2145 35680
rect 1452 35640 1458 35652
rect 2133 35649 2145 35652
rect 2179 35649 2191 35683
rect 19150 35680 19156 35692
rect 19111 35652 19156 35680
rect 2133 35643 2191 35649
rect 19150 35640 19156 35652
rect 19208 35640 19214 35692
rect 19521 35683 19579 35689
rect 19521 35649 19533 35683
rect 19567 35680 19579 35683
rect 19978 35680 19984 35692
rect 19567 35652 19984 35680
rect 19567 35649 19579 35652
rect 19521 35643 19579 35649
rect 19978 35640 19984 35652
rect 20036 35640 20042 35692
rect 20714 35680 20720 35692
rect 20675 35652 20720 35680
rect 20714 35640 20720 35652
rect 20772 35640 20778 35692
rect 21008 35689 21036 35720
rect 20993 35683 21051 35689
rect 20993 35649 21005 35683
rect 21039 35649 21051 35683
rect 20993 35643 21051 35649
rect 21821 35683 21879 35689
rect 21821 35649 21833 35683
rect 21867 35649 21879 35683
rect 21821 35643 21879 35649
rect 22465 35683 22523 35689
rect 22465 35649 22477 35683
rect 22511 35649 22523 35683
rect 22646 35680 22652 35692
rect 22607 35652 22652 35680
rect 22465 35643 22523 35649
rect 19061 35615 19119 35621
rect 9646 35584 17908 35612
rect 8018 35504 8024 35556
rect 8076 35544 8082 35556
rect 9646 35544 9674 35584
rect 8076 35516 9674 35544
rect 17880 35544 17908 35584
rect 19061 35581 19073 35615
rect 19107 35612 19119 35615
rect 20346 35612 20352 35624
rect 19107 35584 20352 35612
rect 19107 35581 19119 35584
rect 19061 35575 19119 35581
rect 20346 35572 20352 35584
rect 20404 35572 20410 35624
rect 20898 35612 20904 35624
rect 20859 35584 20904 35612
rect 20898 35572 20904 35584
rect 20956 35572 20962 35624
rect 21177 35547 21235 35553
rect 17880 35516 19564 35544
rect 8076 35504 8082 35516
rect 1670 35436 1676 35488
rect 1728 35476 1734 35488
rect 14458 35476 14464 35488
rect 1728 35448 14464 35476
rect 1728 35436 1734 35448
rect 14458 35436 14464 35448
rect 14516 35436 14522 35488
rect 19536 35485 19564 35516
rect 21177 35513 21189 35547
rect 21223 35544 21235 35547
rect 21836 35544 21864 35643
rect 22480 35612 22508 35643
rect 22646 35640 22652 35652
rect 22704 35640 22710 35692
rect 23032 35689 23060 35788
rect 23201 35785 23213 35819
rect 23247 35816 23259 35819
rect 36170 35816 36176 35828
rect 23247 35788 36176 35816
rect 23247 35785 23259 35788
rect 23201 35779 23259 35785
rect 36170 35776 36176 35788
rect 36228 35776 36234 35828
rect 36354 35816 36360 35828
rect 36315 35788 36360 35816
rect 36354 35776 36360 35788
rect 36412 35776 36418 35828
rect 37918 35776 37924 35828
rect 37976 35816 37982 35828
rect 38381 35819 38439 35825
rect 38381 35816 38393 35819
rect 37976 35788 38393 35816
rect 37976 35776 37982 35788
rect 38381 35785 38393 35788
rect 38427 35785 38439 35819
rect 67358 35816 67364 35828
rect 38381 35779 38439 35785
rect 41386 35788 67364 35816
rect 25314 35748 25320 35760
rect 24228 35720 25320 35748
rect 24228 35689 24256 35720
rect 25314 35708 25320 35720
rect 25372 35708 25378 35760
rect 28896 35751 28954 35757
rect 28896 35717 28908 35751
rect 28942 35748 28954 35751
rect 29546 35748 29552 35760
rect 28942 35720 29552 35748
rect 28942 35717 28954 35720
rect 28896 35711 28954 35717
rect 29546 35708 29552 35720
rect 29604 35708 29610 35760
rect 32306 35748 32312 35760
rect 31312 35720 32312 35748
rect 24486 35689 24492 35692
rect 23017 35683 23075 35689
rect 23017 35649 23029 35683
rect 23063 35649 23075 35683
rect 23017 35643 23075 35649
rect 24213 35683 24271 35689
rect 24213 35649 24225 35683
rect 24259 35649 24271 35683
rect 24213 35643 24271 35649
rect 24480 35643 24492 35689
rect 24544 35680 24550 35692
rect 27157 35683 27215 35689
rect 24544 35652 24580 35680
rect 24486 35640 24492 35643
rect 24544 35640 24550 35652
rect 27157 35649 27169 35683
rect 27203 35680 27215 35683
rect 27430 35680 27436 35692
rect 27203 35652 27436 35680
rect 27203 35649 27215 35652
rect 27157 35643 27215 35649
rect 27430 35640 27436 35652
rect 27488 35640 27494 35692
rect 28629 35683 28687 35689
rect 28629 35649 28641 35683
rect 28675 35680 28687 35683
rect 28718 35680 28724 35692
rect 28675 35652 28724 35680
rect 28675 35649 28687 35652
rect 28629 35643 28687 35649
rect 28718 35640 28724 35652
rect 28776 35640 28782 35692
rect 30469 35683 30527 35689
rect 30469 35649 30481 35683
rect 30515 35680 30527 35683
rect 30742 35680 30748 35692
rect 30515 35652 30748 35680
rect 30515 35649 30527 35652
rect 30469 35643 30527 35649
rect 30742 35640 30748 35652
rect 30800 35640 30806 35692
rect 31312 35689 31340 35720
rect 32306 35708 32312 35720
rect 32364 35708 32370 35760
rect 41386 35748 41414 35788
rect 67358 35776 67364 35788
rect 67416 35776 67422 35828
rect 42426 35748 42432 35760
rect 35084 35720 41414 35748
rect 42387 35720 42432 35748
rect 31297 35683 31355 35689
rect 31297 35649 31309 35683
rect 31343 35649 31355 35683
rect 31297 35643 31355 35649
rect 31386 35640 31392 35692
rect 31444 35680 31450 35692
rect 32398 35680 32404 35692
rect 31444 35652 31489 35680
rect 31726 35652 32404 35680
rect 31444 35640 31450 35652
rect 22554 35612 22560 35624
rect 22480 35584 22560 35612
rect 22554 35572 22560 35584
rect 22612 35572 22618 35624
rect 31726 35612 31754 35652
rect 32398 35640 32404 35652
rect 32456 35640 32462 35692
rect 33321 35683 33379 35689
rect 33321 35649 33333 35683
rect 33367 35680 33379 35683
rect 33410 35680 33416 35692
rect 33367 35652 33416 35680
rect 33367 35649 33379 35652
rect 33321 35643 33379 35649
rect 33410 35640 33416 35652
rect 33468 35640 33474 35692
rect 30668 35584 31754 35612
rect 30668 35553 30696 35584
rect 30653 35547 30711 35553
rect 21223 35516 21864 35544
rect 25516 35516 27108 35544
rect 21223 35513 21235 35516
rect 21177 35507 21235 35513
rect 19521 35479 19579 35485
rect 19521 35445 19533 35479
rect 19567 35445 19579 35479
rect 19521 35439 19579 35445
rect 20441 35479 20499 35485
rect 20441 35445 20453 35479
rect 20487 35476 20499 35479
rect 20993 35479 21051 35485
rect 20993 35476 21005 35479
rect 20487 35448 21005 35476
rect 20487 35445 20499 35448
rect 20441 35439 20499 35445
rect 20993 35445 21005 35448
rect 21039 35476 21051 35479
rect 25516 35476 25544 35516
rect 21039 35448 25544 35476
rect 25593 35479 25651 35485
rect 21039 35445 21051 35448
rect 20993 35439 21051 35445
rect 25593 35445 25605 35479
rect 25639 35476 25651 35479
rect 25682 35476 25688 35488
rect 25639 35448 25688 35476
rect 25639 35445 25651 35448
rect 25593 35439 25651 35445
rect 25682 35436 25688 35448
rect 25740 35436 25746 35488
rect 26970 35476 26976 35488
rect 26931 35448 26976 35476
rect 26970 35436 26976 35448
rect 27028 35436 27034 35488
rect 27080 35476 27108 35516
rect 29564 35516 30144 35544
rect 29564 35476 29592 35516
rect 30006 35476 30012 35488
rect 27080 35448 29592 35476
rect 29967 35448 30012 35476
rect 30006 35436 30012 35448
rect 30064 35436 30070 35488
rect 30116 35476 30144 35516
rect 30653 35513 30665 35547
rect 30699 35513 30711 35547
rect 35084 35544 35112 35720
rect 42426 35708 42432 35720
rect 42484 35708 42490 35760
rect 42794 35748 42800 35760
rect 42755 35720 42800 35748
rect 42794 35708 42800 35720
rect 42852 35708 42858 35760
rect 46937 35751 46995 35757
rect 46937 35717 46949 35751
rect 46983 35748 46995 35751
rect 48133 35751 48191 35757
rect 48133 35748 48145 35751
rect 46983 35720 48145 35748
rect 46983 35717 46995 35720
rect 46937 35711 46995 35717
rect 48133 35717 48145 35720
rect 48179 35717 48191 35751
rect 66898 35748 66904 35760
rect 48133 35711 48191 35717
rect 65812 35720 66904 35748
rect 35161 35683 35219 35689
rect 35161 35649 35173 35683
rect 35207 35649 35219 35683
rect 35618 35680 35624 35692
rect 35579 35652 35624 35680
rect 35161 35643 35219 35649
rect 35176 35612 35204 35643
rect 35618 35640 35624 35652
rect 35676 35640 35682 35692
rect 36538 35680 36544 35692
rect 36499 35652 36544 35680
rect 36538 35640 36544 35652
rect 36596 35640 36602 35692
rect 37274 35640 37280 35692
rect 37332 35680 37338 35692
rect 38010 35680 38016 35692
rect 37332 35652 38016 35680
rect 37332 35640 37338 35652
rect 38010 35640 38016 35652
rect 38068 35680 38074 35692
rect 38197 35683 38255 35689
rect 38197 35680 38209 35683
rect 38068 35652 38209 35680
rect 38068 35640 38074 35652
rect 38197 35649 38209 35652
rect 38243 35649 38255 35683
rect 39206 35680 39212 35692
rect 39167 35652 39212 35680
rect 38197 35643 38255 35649
rect 39206 35640 39212 35652
rect 39264 35640 39270 35692
rect 39301 35683 39359 35689
rect 39301 35649 39313 35683
rect 39347 35680 39359 35683
rect 40310 35680 40316 35692
rect 39347 35652 40316 35680
rect 39347 35649 39359 35652
rect 39301 35643 39359 35649
rect 40310 35640 40316 35652
rect 40368 35640 40374 35692
rect 40764 35683 40822 35689
rect 40764 35649 40776 35683
rect 40810 35680 40822 35683
rect 41598 35680 41604 35692
rect 40810 35652 41604 35680
rect 40810 35649 40822 35652
rect 40764 35643 40822 35649
rect 41598 35640 41604 35652
rect 41656 35640 41662 35692
rect 42613 35683 42671 35689
rect 42613 35649 42625 35683
rect 42659 35649 42671 35683
rect 42613 35643 42671 35649
rect 43708 35683 43766 35689
rect 43708 35649 43720 35683
rect 43754 35680 43766 35683
rect 43990 35680 43996 35692
rect 43754 35652 43996 35680
rect 43754 35649 43766 35652
rect 43708 35643 43766 35649
rect 35986 35612 35992 35624
rect 35176 35584 35992 35612
rect 35986 35572 35992 35584
rect 36044 35572 36050 35624
rect 40494 35612 40500 35624
rect 40455 35584 40500 35612
rect 40494 35572 40500 35584
rect 40552 35572 40558 35624
rect 42628 35612 42656 35643
rect 43990 35640 43996 35652
rect 44048 35640 44054 35692
rect 46842 35680 46848 35692
rect 46803 35652 46848 35680
rect 46842 35640 46848 35652
rect 46900 35640 46906 35692
rect 47854 35640 47860 35692
rect 47912 35680 47918 35692
rect 65812 35689 65840 35720
rect 66898 35708 66904 35720
rect 66956 35708 66962 35760
rect 47949 35683 48007 35689
rect 47949 35680 47961 35683
rect 47912 35652 47961 35680
rect 47912 35640 47918 35652
rect 47949 35649 47961 35652
rect 47995 35649 48007 35683
rect 47949 35643 48007 35649
rect 65797 35683 65855 35689
rect 65797 35649 65809 35683
rect 65843 35649 65855 35683
rect 65797 35643 65855 35649
rect 42794 35612 42800 35624
rect 41892 35584 42800 35612
rect 30653 35507 30711 35513
rect 30760 35516 35112 35544
rect 30760 35476 30788 35516
rect 35342 35504 35348 35556
rect 35400 35544 35406 35556
rect 41892 35553 41920 35584
rect 42794 35572 42800 35584
rect 42852 35572 42858 35624
rect 43438 35612 43444 35624
rect 43399 35584 43444 35612
rect 43438 35572 43444 35584
rect 43496 35572 43502 35624
rect 49602 35612 49608 35624
rect 49563 35584 49608 35612
rect 49602 35572 49608 35584
rect 49660 35572 49666 35624
rect 65978 35612 65984 35624
rect 65939 35584 65984 35612
rect 65978 35572 65984 35584
rect 66036 35572 66042 35624
rect 67542 35612 67548 35624
rect 67503 35584 67548 35612
rect 67542 35572 67548 35584
rect 67600 35572 67606 35624
rect 35621 35547 35679 35553
rect 35621 35544 35633 35547
rect 35400 35516 35633 35544
rect 35400 35504 35406 35516
rect 35621 35513 35633 35516
rect 35667 35513 35679 35547
rect 35621 35507 35679 35513
rect 41877 35547 41935 35553
rect 41877 35513 41889 35547
rect 41923 35513 41935 35547
rect 44818 35544 44824 35556
rect 44779 35516 44824 35544
rect 41877 35507 41935 35513
rect 44818 35504 44824 35516
rect 44876 35504 44882 35556
rect 30116 35448 30788 35476
rect 31478 35436 31484 35488
rect 31536 35476 31542 35488
rect 31573 35479 31631 35485
rect 31573 35476 31585 35479
rect 31536 35448 31585 35476
rect 31536 35436 31542 35448
rect 31573 35445 31585 35448
rect 31619 35445 31631 35479
rect 32582 35476 32588 35488
rect 32543 35448 32588 35476
rect 31573 35439 31631 35445
rect 32582 35436 32588 35448
rect 32640 35436 32646 35488
rect 33134 35476 33140 35488
rect 33095 35448 33140 35476
rect 33134 35436 33140 35448
rect 33192 35436 33198 35488
rect 34977 35479 35035 35485
rect 34977 35445 34989 35479
rect 35023 35476 35035 35479
rect 35434 35476 35440 35488
rect 35023 35448 35440 35476
rect 35023 35445 35035 35448
rect 34977 35439 35035 35445
rect 35434 35436 35440 35448
rect 35492 35436 35498 35488
rect 35526 35436 35532 35488
rect 35584 35476 35590 35488
rect 35894 35476 35900 35488
rect 35584 35448 35900 35476
rect 35584 35436 35590 35448
rect 35894 35436 35900 35448
rect 35952 35436 35958 35488
rect 39114 35436 39120 35488
rect 39172 35476 39178 35488
rect 39485 35479 39543 35485
rect 39485 35476 39497 35479
rect 39172 35448 39497 35476
rect 39172 35436 39178 35448
rect 39485 35445 39497 35448
rect 39531 35445 39543 35479
rect 39485 35439 39543 35445
rect 1104 35386 68816 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 68816 35386
rect 1104 35312 68816 35334
rect 20070 35232 20076 35284
rect 20128 35272 20134 35284
rect 20165 35275 20223 35281
rect 20165 35272 20177 35275
rect 20128 35244 20177 35272
rect 20128 35232 20134 35244
rect 20165 35241 20177 35244
rect 20211 35241 20223 35275
rect 20165 35235 20223 35241
rect 20625 35275 20683 35281
rect 20625 35241 20637 35275
rect 20671 35272 20683 35275
rect 21726 35272 21732 35284
rect 20671 35244 21732 35272
rect 20671 35241 20683 35244
rect 20625 35235 20683 35241
rect 20180 35136 20208 35235
rect 21726 35232 21732 35244
rect 21784 35232 21790 35284
rect 22278 35272 22284 35284
rect 22239 35244 22284 35272
rect 22278 35232 22284 35244
rect 22336 35232 22342 35284
rect 23014 35272 23020 35284
rect 22975 35244 23020 35272
rect 23014 35232 23020 35244
rect 23072 35232 23078 35284
rect 25682 35272 25688 35284
rect 24504 35244 25688 35272
rect 20993 35207 21051 35213
rect 20993 35173 21005 35207
rect 21039 35204 21051 35207
rect 22646 35204 22652 35216
rect 21039 35176 22652 35204
rect 21039 35173 21051 35176
rect 20993 35167 21051 35173
rect 22646 35164 22652 35176
rect 22704 35164 22710 35216
rect 24504 35145 24532 35244
rect 25682 35232 25688 35244
rect 25740 35272 25746 35284
rect 29733 35275 29791 35281
rect 25740 35244 27936 35272
rect 25740 35232 25746 35244
rect 26697 35207 26755 35213
rect 26697 35173 26709 35207
rect 26743 35204 26755 35207
rect 26743 35176 27200 35204
rect 26743 35173 26755 35176
rect 26697 35167 26755 35173
rect 20625 35139 20683 35145
rect 20625 35136 20637 35139
rect 20180 35108 20637 35136
rect 20625 35105 20637 35108
rect 20671 35105 20683 35139
rect 20625 35099 20683 35105
rect 24489 35139 24547 35145
rect 24489 35105 24501 35139
rect 24535 35105 24547 35139
rect 24489 35099 24547 35105
rect 27062 35096 27068 35148
rect 27120 35136 27126 35148
rect 27172 35145 27200 35176
rect 27706 35164 27712 35216
rect 27764 35204 27770 35216
rect 27801 35207 27859 35213
rect 27801 35204 27813 35207
rect 27764 35176 27813 35204
rect 27764 35164 27770 35176
rect 27801 35173 27813 35176
rect 27847 35173 27859 35207
rect 27801 35167 27859 35173
rect 27157 35139 27215 35145
rect 27157 35136 27169 35139
rect 27120 35108 27169 35136
rect 27120 35096 27126 35108
rect 27157 35105 27169 35108
rect 27203 35105 27215 35139
rect 27157 35099 27215 35105
rect 27341 35139 27399 35145
rect 27341 35105 27353 35139
rect 27387 35105 27399 35139
rect 27908 35136 27936 35244
rect 29733 35241 29745 35275
rect 29779 35241 29791 35275
rect 29914 35272 29920 35284
rect 29875 35244 29920 35272
rect 29733 35235 29791 35241
rect 29748 35204 29776 35235
rect 29914 35232 29920 35244
rect 29972 35232 29978 35284
rect 31294 35272 31300 35284
rect 31255 35244 31300 35272
rect 31294 35232 31300 35244
rect 31352 35232 31358 35284
rect 31570 35232 31576 35284
rect 31628 35272 31634 35284
rect 36541 35275 36599 35281
rect 31628 35244 35480 35272
rect 31628 35232 31634 35244
rect 30466 35204 30472 35216
rect 29748 35176 30472 35204
rect 30466 35164 30472 35176
rect 30524 35164 30530 35216
rect 34514 35164 34520 35216
rect 34572 35204 34578 35216
rect 35345 35207 35403 35213
rect 35345 35204 35357 35207
rect 34572 35176 35357 35204
rect 34572 35164 34578 35176
rect 35345 35173 35357 35176
rect 35391 35173 35403 35207
rect 35345 35167 35403 35173
rect 28194 35139 28252 35145
rect 28194 35136 28206 35139
rect 27908 35108 28206 35136
rect 27341 35099 27399 35105
rect 28194 35105 28206 35108
rect 28240 35105 28252 35139
rect 32582 35136 32588 35148
rect 32543 35108 32588 35136
rect 28194 35099 28252 35105
rect 20806 35068 20812 35080
rect 20767 35040 20812 35068
rect 20806 35028 20812 35040
rect 20864 35028 20870 35080
rect 22370 35068 22376 35080
rect 22331 35040 22376 35068
rect 22370 35028 22376 35040
rect 22428 35028 22434 35080
rect 23201 35071 23259 35077
rect 23201 35037 23213 35071
rect 23247 35068 23259 35071
rect 23750 35068 23756 35080
rect 23247 35040 23756 35068
rect 23247 35037 23259 35040
rect 23201 35031 23259 35037
rect 23750 35028 23756 35040
rect 23808 35028 23814 35080
rect 24673 35071 24731 35077
rect 24673 35037 24685 35071
rect 24719 35037 24731 35071
rect 25314 35068 25320 35080
rect 25275 35040 25320 35068
rect 24673 35031 24731 35037
rect 20530 35000 20536 35012
rect 20491 34972 20536 35000
rect 20530 34960 20536 34972
rect 20588 34960 20594 35012
rect 24688 35000 24716 35031
rect 25314 35028 25320 35040
rect 25372 35028 25378 35080
rect 25584 35071 25642 35077
rect 25584 35037 25596 35071
rect 25630 35068 25642 35071
rect 26970 35068 26976 35080
rect 25630 35040 26976 35068
rect 25630 35037 25642 35040
rect 25584 35031 25642 35037
rect 26970 35028 26976 35040
rect 27028 35028 27034 35080
rect 25498 35000 25504 35012
rect 24688 34972 25504 35000
rect 25498 34960 25504 34972
rect 25556 34960 25562 35012
rect 24854 34932 24860 34944
rect 24815 34904 24860 34932
rect 24854 34892 24860 34904
rect 24912 34892 24918 34944
rect 27356 34932 27384 35099
rect 32582 35096 32588 35108
rect 32640 35096 32646 35148
rect 34885 35139 34943 35145
rect 34885 35105 34897 35139
rect 34931 35136 34943 35139
rect 35250 35136 35256 35148
rect 34931 35108 35256 35136
rect 34931 35105 34943 35108
rect 34885 35099 34943 35105
rect 35250 35096 35256 35108
rect 35308 35096 35314 35148
rect 35452 35136 35480 35244
rect 36541 35241 36553 35275
rect 36587 35272 36599 35275
rect 37366 35272 37372 35284
rect 36587 35244 37372 35272
rect 36587 35241 36599 35244
rect 36541 35235 36599 35241
rect 37366 35232 37372 35244
rect 37424 35232 37430 35284
rect 38930 35272 38936 35284
rect 38891 35244 38936 35272
rect 38930 35232 38936 35244
rect 38988 35232 38994 35284
rect 43438 35232 43444 35284
rect 43496 35272 43502 35284
rect 43625 35275 43683 35281
rect 43625 35272 43637 35275
rect 43496 35244 43637 35272
rect 43496 35232 43502 35244
rect 43625 35241 43637 35244
rect 43671 35241 43683 35275
rect 43625 35235 43683 35241
rect 65978 35232 65984 35284
rect 66036 35272 66042 35284
rect 67545 35275 67603 35281
rect 67545 35272 67557 35275
rect 66036 35244 67557 35272
rect 66036 35232 66042 35244
rect 67545 35241 67557 35244
rect 67591 35241 67603 35275
rect 67545 35235 67603 35241
rect 45646 35204 45652 35216
rect 40144 35176 41414 35204
rect 45607 35176 45652 35204
rect 40144 35148 40172 35176
rect 35738 35139 35796 35145
rect 35738 35136 35750 35139
rect 35452 35108 35750 35136
rect 35738 35105 35750 35108
rect 35784 35105 35796 35139
rect 35894 35136 35900 35148
rect 35855 35108 35900 35136
rect 35738 35099 35796 35105
rect 35894 35096 35900 35108
rect 35952 35096 35958 35148
rect 40126 35136 40132 35148
rect 40087 35108 40132 35136
rect 40126 35096 40132 35108
rect 40184 35096 40190 35148
rect 40310 35096 40316 35148
rect 40368 35136 40374 35148
rect 40405 35139 40463 35145
rect 40405 35136 40417 35139
rect 40368 35108 40417 35136
rect 40368 35096 40374 35108
rect 40405 35105 40417 35108
rect 40451 35105 40463 35139
rect 41386 35136 41414 35176
rect 45646 35164 45652 35176
rect 45704 35164 45710 35216
rect 41509 35139 41567 35145
rect 41509 35136 41521 35139
rect 41386 35108 41521 35136
rect 40405 35099 40463 35105
rect 41509 35105 41521 35108
rect 41555 35105 41567 35139
rect 42794 35136 42800 35148
rect 42755 35108 42800 35136
rect 41509 35099 41567 35105
rect 42794 35096 42800 35108
rect 42852 35096 42858 35148
rect 49234 35136 49240 35148
rect 49195 35108 49240 35136
rect 49234 35096 49240 35108
rect 49292 35096 49298 35148
rect 28074 35028 28080 35080
rect 28132 35068 28138 35080
rect 28350 35068 28356 35080
rect 28132 35040 28177 35068
rect 28311 35040 28356 35068
rect 28132 35028 28138 35040
rect 28350 35028 28356 35040
rect 28408 35028 28414 35080
rect 28997 35071 29055 35077
rect 28997 35037 29009 35071
rect 29043 35068 29055 35071
rect 30561 35071 30619 35077
rect 29043 35040 30328 35068
rect 29043 35037 29055 35040
rect 28997 35031 29055 35037
rect 29549 35003 29607 35009
rect 29549 34969 29561 35003
rect 29595 35000 29607 35003
rect 30006 35000 30012 35012
rect 29595 34972 30012 35000
rect 29595 34969 29607 34972
rect 29549 34963 29607 34969
rect 29564 34932 29592 34963
rect 30006 34960 30012 34972
rect 30064 34960 30070 35012
rect 30300 35000 30328 35040
rect 30561 35037 30573 35071
rect 30607 35068 30619 35071
rect 30834 35068 30840 35080
rect 30607 35040 30840 35068
rect 30607 35037 30619 35040
rect 30561 35031 30619 35037
rect 30834 35028 30840 35040
rect 30892 35028 30898 35080
rect 31478 35068 31484 35080
rect 31439 35040 31484 35068
rect 31478 35028 31484 35040
rect 31536 35028 31542 35080
rect 32852 35071 32910 35077
rect 32852 35037 32864 35071
rect 32898 35068 32910 35071
rect 33134 35068 33140 35080
rect 32898 35040 33140 35068
rect 32898 35037 32910 35040
rect 32852 35031 32910 35037
rect 33134 35028 33140 35040
rect 33192 35028 33198 35080
rect 33962 35028 33968 35080
rect 34020 35068 34026 35080
rect 34701 35071 34759 35077
rect 34701 35068 34713 35071
rect 34020 35040 34713 35068
rect 34020 35028 34026 35040
rect 34701 35037 34713 35040
rect 34747 35037 34759 35071
rect 34701 35031 34759 35037
rect 35618 35028 35624 35080
rect 35676 35068 35682 35080
rect 38473 35071 38531 35077
rect 35676 35040 35721 35068
rect 35676 35028 35682 35040
rect 38473 35037 38485 35071
rect 38519 35068 38531 35071
rect 38930 35068 38936 35080
rect 38519 35040 38936 35068
rect 38519 35037 38531 35040
rect 38473 35031 38531 35037
rect 38930 35028 38936 35040
rect 38988 35028 38994 35080
rect 39114 35068 39120 35080
rect 39075 35040 39120 35068
rect 39114 35028 39120 35040
rect 39172 35028 39178 35080
rect 41785 35071 41843 35077
rect 41785 35037 41797 35071
rect 41831 35068 41843 35071
rect 42978 35068 42984 35080
rect 41831 35040 42984 35068
rect 41831 35037 41843 35040
rect 41785 35031 41843 35037
rect 42978 35028 42984 35040
rect 43036 35028 43042 35080
rect 43625 35071 43683 35077
rect 43625 35037 43637 35071
rect 43671 35037 43683 35071
rect 43625 35031 43683 35037
rect 37185 35003 37243 35009
rect 37185 35000 37197 35003
rect 30300 34972 34468 35000
rect 27356 34904 29592 34932
rect 29730 34892 29736 34944
rect 29788 34941 29794 34944
rect 29788 34935 29807 34941
rect 29795 34901 29807 34935
rect 29788 34895 29807 34901
rect 29788 34892 29794 34895
rect 30190 34892 30196 34944
rect 30248 34932 30254 34944
rect 30561 34935 30619 34941
rect 30561 34932 30573 34935
rect 30248 34904 30573 34932
rect 30248 34892 30254 34904
rect 30561 34901 30573 34904
rect 30607 34901 30619 34935
rect 33962 34932 33968 34944
rect 33923 34904 33968 34932
rect 30561 34895 30619 34901
rect 33962 34892 33968 34904
rect 34020 34892 34026 34944
rect 34440 34932 34468 34972
rect 36372 34972 37197 35000
rect 36372 34932 36400 34972
rect 37185 34969 37197 34972
rect 37231 34969 37243 35003
rect 37185 34963 37243 34969
rect 37369 35003 37427 35009
rect 37369 34969 37381 35003
rect 37415 35000 37427 35003
rect 37458 35000 37464 35012
rect 37415 34972 37464 35000
rect 37415 34969 37427 34972
rect 37369 34963 37427 34969
rect 37458 34960 37464 34972
rect 37516 34960 37522 35012
rect 40954 34960 40960 35012
rect 41012 35000 41018 35012
rect 43640 35000 43668 35031
rect 44266 35028 44272 35080
rect 44324 35068 44330 35080
rect 45278 35068 45284 35080
rect 44324 35040 45284 35068
rect 44324 35028 44330 35040
rect 45278 35028 45284 35040
rect 45336 35068 45342 35080
rect 45465 35071 45523 35077
rect 45465 35068 45477 35071
rect 45336 35040 45477 35068
rect 45336 35028 45342 35040
rect 45465 35037 45477 35040
rect 45511 35037 45523 35071
rect 47486 35068 47492 35080
rect 47447 35040 47492 35068
rect 45465 35031 45523 35037
rect 47486 35028 47492 35040
rect 47544 35028 47550 35080
rect 67450 35068 67456 35080
rect 67411 35040 67456 35068
rect 67450 35028 67456 35040
rect 67508 35028 67514 35080
rect 47670 35000 47676 35012
rect 41012 34972 43668 35000
rect 47631 34972 47676 35000
rect 41012 34960 41018 34972
rect 47670 34960 47676 34972
rect 47728 34960 47734 35012
rect 34440 34904 36400 34932
rect 37553 34935 37611 34941
rect 37553 34901 37565 34935
rect 37599 34932 37611 34935
rect 38010 34932 38016 34944
rect 37599 34904 38016 34932
rect 37599 34901 37611 34904
rect 37553 34895 37611 34901
rect 38010 34892 38016 34904
rect 38068 34892 38074 34944
rect 38102 34892 38108 34944
rect 38160 34932 38166 34944
rect 38289 34935 38347 34941
rect 38289 34932 38301 34935
rect 38160 34904 38301 34932
rect 38160 34892 38166 34904
rect 38289 34901 38301 34904
rect 38335 34901 38347 34935
rect 38289 34895 38347 34901
rect 41782 34892 41788 34944
rect 41840 34932 41846 34944
rect 43165 34935 43223 34941
rect 43165 34932 43177 34935
rect 41840 34904 43177 34932
rect 41840 34892 41846 34904
rect 43165 34901 43177 34904
rect 43211 34901 43223 34935
rect 43165 34895 43223 34901
rect 1104 34842 68816 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 68816 34842
rect 1104 34768 68816 34790
rect 24486 34688 24492 34740
rect 24544 34728 24550 34740
rect 24673 34731 24731 34737
rect 24673 34728 24685 34731
rect 24544 34700 24685 34728
rect 24544 34688 24550 34700
rect 24673 34697 24685 34700
rect 24719 34697 24731 34731
rect 24673 34691 24731 34697
rect 25314 34688 25320 34740
rect 25372 34728 25378 34740
rect 25961 34731 26019 34737
rect 25961 34728 25973 34731
rect 25372 34700 25973 34728
rect 25372 34688 25378 34700
rect 25961 34697 25973 34700
rect 26007 34697 26019 34731
rect 27430 34728 27436 34740
rect 27391 34700 27436 34728
rect 25961 34691 26019 34697
rect 27430 34688 27436 34700
rect 27488 34688 27494 34740
rect 31570 34728 31576 34740
rect 31531 34700 31576 34728
rect 31570 34688 31576 34700
rect 31628 34688 31634 34740
rect 32125 34731 32183 34737
rect 32125 34728 32137 34731
rect 31726 34700 32137 34728
rect 27062 34660 27068 34672
rect 27023 34632 27068 34660
rect 27062 34620 27068 34632
rect 27120 34620 27126 34672
rect 27281 34663 27339 34669
rect 27281 34629 27293 34663
rect 27327 34660 27339 34663
rect 28810 34660 28816 34672
rect 27327 34632 28816 34660
rect 27327 34629 27339 34632
rect 27281 34623 27339 34629
rect 28810 34620 28816 34632
rect 28868 34620 28874 34672
rect 30460 34663 30518 34669
rect 30460 34629 30472 34663
rect 30506 34660 30518 34663
rect 31726 34660 31754 34700
rect 32125 34697 32137 34700
rect 32171 34697 32183 34731
rect 33410 34728 33416 34740
rect 33371 34700 33416 34728
rect 32125 34691 32183 34697
rect 33410 34688 33416 34700
rect 33468 34688 33474 34740
rect 35250 34688 35256 34740
rect 35308 34728 35314 34740
rect 36725 34731 36783 34737
rect 36725 34728 36737 34731
rect 35308 34700 36737 34728
rect 35308 34688 35314 34700
rect 36725 34697 36737 34700
rect 36771 34697 36783 34731
rect 36725 34691 36783 34697
rect 38933 34731 38991 34737
rect 38933 34697 38945 34731
rect 38979 34728 38991 34731
rect 40218 34728 40224 34740
rect 38979 34700 40224 34728
rect 38979 34697 38991 34700
rect 38933 34691 38991 34697
rect 40218 34688 40224 34700
rect 40276 34688 40282 34740
rect 40494 34688 40500 34740
rect 40552 34728 40558 34740
rect 40957 34731 41015 34737
rect 40957 34728 40969 34731
rect 40552 34700 40969 34728
rect 40552 34688 40558 34700
rect 40957 34697 40969 34700
rect 41003 34697 41015 34731
rect 41598 34728 41604 34740
rect 41559 34700 41604 34728
rect 40957 34691 41015 34697
rect 41598 34688 41604 34700
rect 41656 34688 41662 34740
rect 43990 34728 43996 34740
rect 43951 34700 43996 34728
rect 43990 34688 43996 34700
rect 44048 34688 44054 34740
rect 45370 34688 45376 34740
rect 45428 34728 45434 34740
rect 46845 34731 46903 34737
rect 46845 34728 46857 34731
rect 45428 34700 46857 34728
rect 45428 34688 45434 34700
rect 46845 34697 46857 34700
rect 46891 34728 46903 34731
rect 47486 34728 47492 34740
rect 46891 34700 47492 34728
rect 46891 34697 46903 34700
rect 46845 34691 46903 34697
rect 47486 34688 47492 34700
rect 47544 34688 47550 34740
rect 47670 34728 47676 34740
rect 47631 34700 47676 34728
rect 47670 34688 47676 34700
rect 47728 34688 47734 34740
rect 30506 34632 31754 34660
rect 33045 34663 33103 34669
rect 30506 34629 30518 34632
rect 30460 34623 30518 34629
rect 33045 34629 33057 34663
rect 33091 34629 33103 34663
rect 33045 34623 33103 34629
rect 1673 34595 1731 34601
rect 1673 34561 1685 34595
rect 1719 34592 1731 34595
rect 20530 34592 20536 34604
rect 1719 34564 20536 34592
rect 1719 34561 1731 34564
rect 1673 34555 1731 34561
rect 20530 34552 20536 34564
rect 20588 34552 20594 34604
rect 23109 34595 23167 34601
rect 23109 34561 23121 34595
rect 23155 34592 23167 34595
rect 23474 34592 23480 34604
rect 23155 34564 23480 34592
rect 23155 34561 23167 34564
rect 23109 34555 23167 34561
rect 23474 34552 23480 34564
rect 23532 34552 23538 34604
rect 24854 34592 24860 34604
rect 24815 34564 24860 34592
rect 24854 34552 24860 34564
rect 24912 34552 24918 34604
rect 25961 34595 26019 34601
rect 25961 34561 25973 34595
rect 26007 34592 26019 34595
rect 26050 34592 26056 34604
rect 26007 34564 26056 34592
rect 26007 34561 26019 34564
rect 25961 34555 26019 34561
rect 26050 34552 26056 34564
rect 26108 34552 26114 34604
rect 30190 34592 30196 34604
rect 30151 34564 30196 34592
rect 30190 34552 30196 34564
rect 30248 34552 30254 34604
rect 32306 34592 32312 34604
rect 32267 34564 32312 34592
rect 32306 34552 32312 34564
rect 32364 34552 32370 34604
rect 33060 34592 33088 34623
rect 33226 34620 33232 34672
rect 33284 34669 33290 34672
rect 33284 34663 33303 34669
rect 33291 34629 33303 34663
rect 37734 34660 37740 34672
rect 37695 34632 37740 34660
rect 33284 34623 33303 34629
rect 33284 34620 33290 34623
rect 37734 34620 37740 34632
rect 37792 34620 37798 34672
rect 33962 34592 33968 34604
rect 33060 34564 33968 34592
rect 33962 34552 33968 34564
rect 34020 34552 34026 34604
rect 35342 34592 35348 34604
rect 35303 34564 35348 34592
rect 35342 34552 35348 34564
rect 35400 34552 35406 34604
rect 35434 34552 35440 34604
rect 35492 34592 35498 34604
rect 35601 34595 35659 34601
rect 35601 34592 35613 34595
rect 35492 34564 35613 34592
rect 35492 34552 35498 34564
rect 35601 34561 35613 34564
rect 35647 34561 35659 34595
rect 35601 34555 35659 34561
rect 38010 34552 38016 34604
rect 38068 34592 38074 34604
rect 39209 34595 39267 34601
rect 39209 34592 39221 34595
rect 38068 34564 39221 34592
rect 38068 34552 38074 34564
rect 39209 34561 39221 34564
rect 39255 34561 39267 34595
rect 39209 34555 39267 34561
rect 39301 34595 39359 34601
rect 39301 34561 39313 34595
rect 39347 34592 39359 34595
rect 39482 34592 39488 34604
rect 39347 34564 39488 34592
rect 39347 34561 39359 34564
rect 39301 34555 39359 34561
rect 39482 34552 39488 34564
rect 39540 34552 39546 34604
rect 40954 34592 40960 34604
rect 40915 34564 40960 34592
rect 40954 34552 40960 34564
rect 41012 34552 41018 34604
rect 41782 34592 41788 34604
rect 41743 34564 41788 34592
rect 41782 34552 41788 34564
rect 41840 34552 41846 34604
rect 44174 34592 44180 34604
rect 44135 34564 44180 34592
rect 44174 34552 44180 34564
rect 44232 34552 44238 34604
rect 45465 34595 45523 34601
rect 45465 34561 45477 34595
rect 45511 34592 45523 34595
rect 45554 34592 45560 34604
rect 45511 34564 45560 34592
rect 45511 34561 45523 34564
rect 45465 34555 45523 34561
rect 45554 34552 45560 34564
rect 45612 34552 45618 34604
rect 45738 34601 45744 34604
rect 45732 34555 45744 34601
rect 45796 34592 45802 34604
rect 45796 34564 45832 34592
rect 45738 34552 45744 34555
rect 45796 34552 45802 34564
rect 46750 34552 46756 34604
rect 46808 34592 46814 34604
rect 47581 34595 47639 34601
rect 47581 34592 47593 34595
rect 46808 34564 47593 34592
rect 46808 34552 46814 34564
rect 47581 34561 47593 34564
rect 47627 34561 47639 34595
rect 67266 34592 67272 34604
rect 67227 34564 67272 34592
rect 47581 34555 47639 34561
rect 67266 34552 67272 34564
rect 67324 34552 67330 34604
rect 1394 34524 1400 34536
rect 1355 34496 1400 34524
rect 1394 34484 1400 34496
rect 1452 34484 1458 34536
rect 39114 34524 39120 34536
rect 39075 34496 39120 34524
rect 39114 34484 39120 34496
rect 39172 34484 39178 34536
rect 39390 34484 39396 34536
rect 39448 34524 39454 34536
rect 39448 34496 39493 34524
rect 39448 34484 39454 34496
rect 37182 34416 37188 34468
rect 37240 34456 37246 34468
rect 37240 34428 45508 34456
rect 37240 34416 37246 34428
rect 22738 34348 22744 34400
rect 22796 34388 22802 34400
rect 22925 34391 22983 34397
rect 22925 34388 22937 34391
rect 22796 34360 22937 34388
rect 22796 34348 22802 34360
rect 22925 34357 22937 34360
rect 22971 34357 22983 34391
rect 22925 34351 22983 34357
rect 27249 34391 27307 34397
rect 27249 34357 27261 34391
rect 27295 34388 27307 34391
rect 27338 34388 27344 34400
rect 27295 34360 27344 34388
rect 27295 34357 27307 34360
rect 27249 34351 27307 34357
rect 27338 34348 27344 34360
rect 27396 34388 27402 34400
rect 28166 34388 28172 34400
rect 27396 34360 28172 34388
rect 27396 34348 27402 34360
rect 28166 34348 28172 34360
rect 28224 34348 28230 34400
rect 33134 34348 33140 34400
rect 33192 34388 33198 34400
rect 33229 34391 33287 34397
rect 33229 34388 33241 34391
rect 33192 34360 33241 34388
rect 33192 34348 33198 34360
rect 33229 34357 33241 34360
rect 33275 34357 33287 34391
rect 37826 34388 37832 34400
rect 37787 34360 37832 34388
rect 33229 34351 33287 34357
rect 37826 34348 37832 34360
rect 37884 34348 37890 34400
rect 45480 34388 45508 34428
rect 46400 34428 55214 34456
rect 46400 34388 46428 34428
rect 45480 34360 46428 34388
rect 55186 34388 55214 34428
rect 67361 34391 67419 34397
rect 67361 34388 67373 34391
rect 55186 34360 67373 34388
rect 67361 34357 67373 34360
rect 67407 34357 67419 34391
rect 67361 34351 67419 34357
rect 1104 34298 68816 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 68816 34298
rect 1104 34224 68816 34246
rect 23382 34144 23388 34196
rect 23440 34184 23446 34196
rect 23845 34187 23903 34193
rect 23845 34184 23857 34187
rect 23440 34156 23857 34184
rect 23440 34144 23446 34156
rect 23845 34153 23857 34156
rect 23891 34184 23903 34187
rect 28074 34184 28080 34196
rect 23891 34156 28080 34184
rect 23891 34153 23903 34156
rect 23845 34147 23903 34153
rect 28074 34144 28080 34156
rect 28132 34144 28138 34196
rect 28350 34144 28356 34196
rect 28408 34184 28414 34196
rect 28534 34184 28540 34196
rect 28408 34156 28540 34184
rect 28408 34144 28414 34156
rect 28534 34144 28540 34156
rect 28592 34144 28598 34196
rect 30466 34184 30472 34196
rect 30379 34156 30472 34184
rect 30466 34144 30472 34156
rect 30524 34184 30530 34196
rect 30834 34184 30840 34196
rect 30524 34156 30840 34184
rect 30524 34144 30530 34156
rect 30834 34144 30840 34156
rect 30892 34144 30898 34196
rect 31481 34187 31539 34193
rect 31481 34153 31493 34187
rect 31527 34184 31539 34187
rect 32306 34184 32312 34196
rect 31527 34156 32312 34184
rect 31527 34153 31539 34156
rect 31481 34147 31539 34153
rect 32306 34144 32312 34156
rect 32364 34144 32370 34196
rect 35710 34144 35716 34196
rect 35768 34184 35774 34196
rect 35805 34187 35863 34193
rect 35805 34184 35817 34187
rect 35768 34156 35817 34184
rect 35768 34144 35774 34156
rect 35805 34153 35817 34156
rect 35851 34153 35863 34187
rect 35986 34184 35992 34196
rect 35947 34156 35992 34184
rect 35805 34147 35863 34153
rect 35986 34144 35992 34156
rect 36044 34144 36050 34196
rect 45097 34187 45155 34193
rect 45097 34153 45109 34187
rect 45143 34184 45155 34187
rect 45738 34184 45744 34196
rect 45143 34156 45744 34184
rect 45143 34153 45155 34156
rect 45097 34147 45155 34153
rect 45738 34144 45744 34156
rect 45796 34144 45802 34196
rect 33778 34116 33784 34128
rect 29564 34088 33784 34116
rect 22462 33980 22468 33992
rect 22423 33952 22468 33980
rect 22462 33940 22468 33952
rect 22520 33940 22526 33992
rect 22738 33989 22744 33992
rect 22732 33980 22744 33989
rect 22699 33952 22744 33980
rect 22732 33943 22744 33952
rect 22738 33940 22744 33943
rect 22796 33940 22802 33992
rect 24581 33983 24639 33989
rect 24581 33949 24593 33983
rect 24627 33980 24639 33983
rect 24946 33980 24952 33992
rect 24627 33952 24952 33980
rect 24627 33949 24639 33952
rect 24581 33943 24639 33949
rect 24946 33940 24952 33952
rect 25004 33940 25010 33992
rect 25314 33980 25320 33992
rect 25275 33952 25320 33980
rect 25314 33940 25320 33952
rect 25372 33940 25378 33992
rect 28258 33940 28264 33992
rect 28316 33980 28322 33992
rect 28353 33983 28411 33989
rect 28353 33980 28365 33983
rect 28316 33952 28365 33980
rect 28316 33940 28322 33952
rect 28353 33949 28365 33952
rect 28399 33980 28411 33983
rect 28902 33980 28908 33992
rect 28399 33952 28908 33980
rect 28399 33949 28411 33952
rect 28353 33943 28411 33949
rect 28902 33940 28908 33952
rect 28960 33940 28966 33992
rect 29564 33989 29592 34088
rect 33778 34076 33784 34088
rect 33836 34076 33842 34128
rect 42794 34116 42800 34128
rect 42720 34088 42800 34116
rect 31113 34051 31171 34057
rect 31113 34017 31125 34051
rect 31159 34048 31171 34051
rect 31570 34048 31576 34060
rect 31159 34020 31576 34048
rect 31159 34017 31171 34020
rect 31113 34011 31171 34017
rect 31570 34008 31576 34020
rect 31628 34008 31634 34060
rect 40402 34048 40408 34060
rect 40363 34020 40408 34048
rect 40402 34008 40408 34020
rect 40460 34008 40466 34060
rect 42720 34057 42748 34088
rect 42794 34076 42800 34088
rect 42852 34076 42858 34128
rect 42705 34051 42763 34057
rect 42705 34017 42717 34051
rect 42751 34017 42763 34051
rect 42705 34011 42763 34017
rect 42889 34051 42947 34057
rect 42889 34017 42901 34051
rect 42935 34048 42947 34051
rect 43254 34048 43260 34060
rect 42935 34020 43260 34048
rect 42935 34017 42947 34020
rect 42889 34011 42947 34017
rect 43254 34008 43260 34020
rect 43312 34008 43318 34060
rect 44008 34020 45600 34048
rect 29549 33983 29607 33989
rect 29549 33949 29561 33983
rect 29595 33949 29607 33983
rect 29549 33943 29607 33949
rect 29638 33940 29644 33992
rect 29696 33980 29702 33992
rect 30285 33983 30343 33989
rect 30285 33980 30297 33983
rect 29696 33952 30297 33980
rect 29696 33940 29702 33952
rect 30285 33949 30297 33952
rect 30331 33949 30343 33983
rect 30285 33943 30343 33949
rect 31297 33983 31355 33989
rect 31297 33949 31309 33983
rect 31343 33980 31355 33983
rect 31386 33980 31392 33992
rect 31343 33952 31392 33980
rect 31343 33949 31355 33952
rect 31297 33943 31355 33949
rect 31386 33940 31392 33952
rect 31444 33940 31450 33992
rect 37185 33983 37243 33989
rect 37185 33949 37197 33983
rect 37231 33980 37243 33983
rect 37274 33980 37280 33992
rect 37231 33952 37280 33980
rect 37231 33949 37243 33952
rect 37185 33943 37243 33949
rect 37274 33940 37280 33952
rect 37332 33940 37338 33992
rect 38102 33989 38108 33992
rect 37369 33983 37427 33989
rect 37369 33949 37381 33983
rect 37415 33980 37427 33983
rect 37829 33983 37887 33989
rect 37829 33980 37841 33983
rect 37415 33952 37841 33980
rect 37415 33949 37427 33952
rect 37369 33943 37427 33949
rect 37829 33949 37841 33952
rect 37875 33949 37887 33983
rect 38096 33980 38108 33989
rect 38063 33952 38108 33980
rect 37829 33943 37887 33949
rect 38096 33943 38108 33952
rect 38102 33940 38108 33943
rect 38160 33940 38166 33992
rect 40420 33980 40448 34008
rect 40420 33952 41368 33980
rect 41340 33924 41368 33952
rect 42058 33940 42064 33992
rect 42116 33980 42122 33992
rect 42797 33983 42855 33989
rect 42797 33980 42809 33983
rect 42116 33952 42809 33980
rect 42116 33940 42122 33952
rect 42797 33949 42809 33952
rect 42843 33949 42855 33983
rect 42797 33943 42855 33949
rect 42981 33983 43039 33989
rect 42981 33949 42993 33983
rect 43027 33980 43039 33983
rect 43070 33980 43076 33992
rect 43027 33952 43076 33980
rect 43027 33949 43039 33952
rect 42981 33943 43039 33949
rect 43070 33940 43076 33952
rect 43128 33940 43134 33992
rect 43162 33940 43168 33992
rect 43220 33980 43226 33992
rect 43901 33983 43959 33989
rect 43901 33980 43913 33983
rect 43220 33952 43913 33980
rect 43220 33940 43226 33952
rect 43901 33949 43913 33952
rect 43947 33949 43959 33983
rect 43901 33943 43959 33949
rect 29748 33884 31754 33912
rect 24394 33804 24400 33856
rect 24452 33844 24458 33856
rect 24581 33847 24639 33853
rect 24581 33844 24593 33847
rect 24452 33816 24593 33844
rect 24452 33804 24458 33816
rect 24581 33813 24593 33816
rect 24627 33813 24639 33847
rect 25130 33844 25136 33856
rect 25091 33816 25136 33844
rect 24581 33807 24639 33813
rect 25130 33804 25136 33816
rect 25188 33804 25194 33856
rect 29748 33853 29776 33884
rect 29733 33847 29791 33853
rect 29733 33813 29745 33847
rect 29779 33813 29791 33847
rect 31726 33844 31754 33884
rect 35342 33872 35348 33924
rect 35400 33912 35406 33924
rect 35621 33915 35679 33921
rect 35621 33912 35633 33915
rect 35400 33884 35633 33912
rect 35400 33872 35406 33884
rect 35621 33881 35633 33884
rect 35667 33881 35679 33915
rect 35621 33875 35679 33881
rect 40034 33872 40040 33924
rect 40092 33912 40098 33924
rect 40650 33915 40708 33921
rect 40650 33912 40662 33915
rect 40092 33884 40662 33912
rect 40092 33872 40098 33884
rect 40650 33881 40662 33884
rect 40696 33881 40708 33915
rect 40650 33875 40708 33881
rect 41322 33872 41328 33924
rect 41380 33872 41386 33924
rect 44008 33912 44036 34020
rect 45370 33980 45376 33992
rect 45331 33952 45376 33980
rect 45370 33940 45376 33952
rect 45428 33940 45434 33992
rect 45572 33989 45600 34020
rect 45465 33983 45523 33989
rect 45465 33949 45477 33983
rect 45511 33949 45523 33983
rect 45465 33943 45523 33949
rect 45557 33983 45615 33989
rect 45557 33949 45569 33983
rect 45603 33949 45615 33983
rect 45557 33943 45615 33949
rect 42766 33884 44036 33912
rect 34054 33844 34060 33856
rect 31726 33816 34060 33844
rect 29733 33807 29791 33813
rect 34054 33804 34060 33816
rect 34112 33804 34118 33856
rect 35802 33804 35808 33856
rect 35860 33853 35866 33856
rect 35860 33847 35879 33853
rect 35867 33813 35879 33847
rect 35860 33807 35879 33813
rect 35860 33804 35866 33807
rect 39022 33804 39028 33856
rect 39080 33844 39086 33856
rect 39209 33847 39267 33853
rect 39209 33844 39221 33847
rect 39080 33816 39221 33844
rect 39080 33804 39086 33816
rect 39209 33813 39221 33816
rect 39255 33813 39267 33847
rect 39209 33807 39267 33813
rect 41230 33804 41236 33856
rect 41288 33844 41294 33856
rect 41785 33847 41843 33853
rect 41785 33844 41797 33847
rect 41288 33816 41797 33844
rect 41288 33804 41294 33816
rect 41785 33813 41797 33816
rect 41831 33813 41843 33847
rect 41785 33807 41843 33813
rect 42521 33847 42579 33853
rect 42521 33813 42533 33847
rect 42567 33844 42579 33847
rect 42766 33844 42794 33884
rect 44450 33872 44456 33924
rect 44508 33912 44514 33924
rect 45186 33912 45192 33924
rect 44508 33884 45192 33912
rect 44508 33872 44514 33884
rect 45186 33872 45192 33884
rect 45244 33912 45250 33924
rect 45480 33912 45508 33943
rect 45646 33940 45652 33992
rect 45704 33980 45710 33992
rect 45741 33983 45799 33989
rect 45741 33980 45753 33983
rect 45704 33952 45753 33980
rect 45704 33940 45710 33952
rect 45741 33949 45753 33952
rect 45787 33949 45799 33983
rect 45741 33943 45799 33949
rect 45244 33884 45508 33912
rect 45244 33872 45250 33884
rect 43714 33844 43720 33856
rect 42567 33816 42794 33844
rect 43675 33816 43720 33844
rect 42567 33813 42579 33816
rect 42521 33807 42579 33813
rect 43714 33804 43720 33816
rect 43772 33804 43778 33856
rect 1104 33754 68816 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 68816 33754
rect 1104 33680 68816 33702
rect 22462 33600 22468 33652
rect 22520 33640 22526 33652
rect 22557 33643 22615 33649
rect 22557 33640 22569 33643
rect 22520 33612 22569 33640
rect 22520 33600 22526 33612
rect 22557 33609 22569 33612
rect 22603 33609 22615 33643
rect 23474 33640 23480 33652
rect 23435 33612 23480 33640
rect 22557 33603 22615 33609
rect 23474 33600 23480 33612
rect 23532 33600 23538 33652
rect 30098 33640 30104 33652
rect 27540 33612 30104 33640
rect 23382 33572 23388 33584
rect 23216 33544 23388 33572
rect 22370 33504 22376 33516
rect 22331 33476 22376 33504
rect 22370 33464 22376 33476
rect 22428 33464 22434 33516
rect 23216 33513 23244 33544
rect 23382 33532 23388 33544
rect 23440 33532 23446 33584
rect 24664 33575 24722 33581
rect 24664 33541 24676 33575
rect 24710 33572 24722 33575
rect 25130 33572 25136 33584
rect 24710 33544 25136 33572
rect 24710 33541 24722 33544
rect 24664 33535 24722 33541
rect 25130 33532 25136 33544
rect 25188 33532 25194 33584
rect 23201 33507 23259 33513
rect 23201 33473 23213 33507
rect 23247 33473 23259 33507
rect 23201 33467 23259 33473
rect 23293 33507 23351 33513
rect 23293 33473 23305 33507
rect 23339 33504 23351 33507
rect 23566 33504 23572 33516
rect 23339 33476 23572 33504
rect 23339 33473 23351 33476
rect 23293 33467 23351 33473
rect 23566 33464 23572 33476
rect 23624 33464 23630 33516
rect 24394 33504 24400 33516
rect 24355 33476 24400 33504
rect 24394 33464 24400 33476
rect 24452 33464 24458 33516
rect 27540 33513 27568 33612
rect 30098 33600 30104 33612
rect 30156 33600 30162 33652
rect 38473 33643 38531 33649
rect 38473 33609 38485 33643
rect 38519 33640 38531 33643
rect 39114 33640 39120 33652
rect 38519 33612 39120 33640
rect 38519 33609 38531 33612
rect 38473 33603 38531 33609
rect 39114 33600 39120 33612
rect 39172 33600 39178 33652
rect 40034 33640 40040 33652
rect 39995 33612 40040 33640
rect 40034 33600 40040 33612
rect 40092 33600 40098 33652
rect 40310 33640 40316 33652
rect 40144 33612 40316 33640
rect 33226 33581 33232 33584
rect 32953 33575 33011 33581
rect 32953 33541 32965 33575
rect 32999 33541 33011 33575
rect 32953 33535 33011 33541
rect 33169 33575 33232 33581
rect 33169 33541 33181 33575
rect 33215 33541 33232 33575
rect 33169 33535 33232 33541
rect 27525 33507 27583 33513
rect 27525 33473 27537 33507
rect 27571 33473 27583 33507
rect 28534 33504 28540 33516
rect 28495 33476 28540 33504
rect 27525 33467 27583 33473
rect 28534 33464 28540 33476
rect 28592 33464 28598 33516
rect 29641 33507 29699 33513
rect 29641 33473 29653 33507
rect 29687 33473 29699 33507
rect 30466 33504 30472 33516
rect 30427 33476 30472 33504
rect 29641 33467 29699 33473
rect 27341 33439 27399 33445
rect 27341 33405 27353 33439
rect 27387 33405 27399 33439
rect 27341 33399 27399 33405
rect 27356 33368 27384 33399
rect 27706 33396 27712 33448
rect 27764 33436 27770 33448
rect 27985 33439 28043 33445
rect 27985 33436 27997 33439
rect 27764 33408 27997 33436
rect 27764 33396 27770 33408
rect 27985 33405 27997 33408
rect 28031 33405 28043 33439
rect 28258 33436 28264 33448
rect 28219 33408 28264 33436
rect 27985 33399 28043 33405
rect 28258 33396 28264 33408
rect 28316 33396 28322 33448
rect 28350 33396 28356 33448
rect 28408 33445 28414 33448
rect 28408 33439 28436 33445
rect 28424 33405 28436 33439
rect 28408 33399 28436 33405
rect 28408 33396 28414 33399
rect 28902 33396 28908 33448
rect 28960 33436 28966 33448
rect 29656 33436 29684 33467
rect 30466 33464 30472 33476
rect 30524 33464 30530 33516
rect 32968 33504 32996 33535
rect 33226 33532 33232 33535
rect 33284 33532 33290 33584
rect 38105 33575 38163 33581
rect 38105 33541 38117 33575
rect 38151 33572 38163 33575
rect 38838 33572 38844 33584
rect 38151 33544 38844 33572
rect 38151 33541 38163 33544
rect 38105 33535 38163 33541
rect 38838 33532 38844 33544
rect 38896 33532 38902 33584
rect 38930 33532 38936 33584
rect 38988 33572 38994 33584
rect 39301 33575 39359 33581
rect 39301 33572 39313 33575
rect 38988 33544 39313 33572
rect 38988 33532 38994 33544
rect 39301 33541 39313 33544
rect 39347 33541 39359 33575
rect 39301 33535 39359 33541
rect 33778 33504 33784 33516
rect 32968 33476 33784 33504
rect 33778 33464 33784 33476
rect 33836 33464 33842 33516
rect 35621 33507 35679 33513
rect 35621 33473 35633 33507
rect 35667 33504 35679 33507
rect 35710 33504 35716 33516
rect 35667 33476 35716 33504
rect 35667 33473 35679 33476
rect 35621 33467 35679 33473
rect 35710 33464 35716 33476
rect 35768 33464 35774 33516
rect 38289 33507 38347 33513
rect 38289 33473 38301 33507
rect 38335 33504 38347 33507
rect 39022 33504 39028 33516
rect 38335 33476 39028 33504
rect 38335 33473 38347 33476
rect 38289 33467 38347 33473
rect 39022 33464 39028 33476
rect 39080 33464 39086 33516
rect 39117 33507 39175 33513
rect 39117 33473 39129 33507
rect 39163 33504 39175 33507
rect 40034 33504 40040 33516
rect 39163 33476 40040 33504
rect 39163 33473 39175 33476
rect 39117 33467 39175 33473
rect 40034 33464 40040 33476
rect 40092 33504 40098 33516
rect 40144 33504 40172 33612
rect 40310 33600 40316 33612
rect 40368 33600 40374 33652
rect 43162 33640 43168 33652
rect 43123 33612 43168 33640
rect 43162 33600 43168 33612
rect 43220 33600 43226 33652
rect 45005 33643 45063 33649
rect 45005 33640 45017 33643
rect 43272 33612 45017 33640
rect 40218 33532 40224 33584
rect 40276 33572 40282 33584
rect 43272 33572 43300 33612
rect 45005 33609 45017 33612
rect 45051 33609 45063 33643
rect 45005 33603 45063 33609
rect 40276 33544 40540 33572
rect 40276 33532 40282 33544
rect 40512 33513 40540 33544
rect 42904 33544 43300 33572
rect 40313 33507 40371 33513
rect 40313 33504 40325 33507
rect 40092 33476 40172 33504
rect 40236 33476 40325 33504
rect 40092 33464 40098 33476
rect 28960 33408 29684 33436
rect 28960 33396 28966 33408
rect 33042 33396 33048 33448
rect 33100 33436 33106 33448
rect 35345 33439 35403 33445
rect 35345 33436 35357 33439
rect 33100 33408 35357 33436
rect 33100 33396 33106 33408
rect 35345 33405 35357 33408
rect 35391 33436 35403 33439
rect 35434 33436 35440 33448
rect 35391 33408 35440 33436
rect 35391 33405 35403 33408
rect 35345 33399 35403 33405
rect 35434 33396 35440 33408
rect 35492 33396 35498 33448
rect 27614 33368 27620 33380
rect 27356 33340 27620 33368
rect 27614 33328 27620 33340
rect 27672 33328 27678 33380
rect 29181 33371 29239 33377
rect 29181 33337 29193 33371
rect 29227 33368 29239 33371
rect 37366 33368 37372 33380
rect 29227 33340 37372 33368
rect 29227 33337 29239 33340
rect 29181 33331 29239 33337
rect 37366 33328 37372 33340
rect 37424 33328 37430 33380
rect 25774 33300 25780 33312
rect 25687 33272 25780 33300
rect 25774 33260 25780 33272
rect 25832 33300 25838 33312
rect 28350 33300 28356 33312
rect 25832 33272 28356 33300
rect 25832 33260 25838 33272
rect 28350 33260 28356 33272
rect 28408 33260 28414 33312
rect 29822 33300 29828 33312
rect 29783 33272 29828 33300
rect 29822 33260 29828 33272
rect 29880 33260 29886 33312
rect 30558 33300 30564 33312
rect 30519 33272 30564 33300
rect 30558 33260 30564 33272
rect 30616 33260 30622 33312
rect 33134 33300 33140 33312
rect 33095 33272 33140 33300
rect 33134 33260 33140 33272
rect 33192 33260 33198 33312
rect 33318 33300 33324 33312
rect 33279 33272 33324 33300
rect 33318 33260 33324 33272
rect 33376 33260 33382 33312
rect 40236 33300 40264 33476
rect 40313 33473 40325 33476
rect 40359 33473 40371 33507
rect 40313 33467 40371 33473
rect 40405 33507 40463 33513
rect 40405 33473 40417 33507
rect 40451 33473 40463 33507
rect 40405 33467 40463 33473
rect 40497 33507 40555 33513
rect 40497 33473 40509 33507
rect 40543 33473 40555 33507
rect 40678 33504 40684 33516
rect 40639 33476 40684 33504
rect 40497 33467 40555 33473
rect 40420 33436 40448 33467
rect 40678 33464 40684 33476
rect 40736 33464 40742 33516
rect 42794 33464 42800 33516
rect 42852 33504 42858 33516
rect 42904 33513 42932 33544
rect 43714 33532 43720 33584
rect 43772 33572 43778 33584
rect 43870 33575 43928 33581
rect 43870 33572 43882 33575
rect 43772 33544 43882 33572
rect 43772 33532 43778 33544
rect 43870 33541 43882 33544
rect 43916 33541 43928 33575
rect 43870 33535 43928 33541
rect 42889 33507 42947 33513
rect 42889 33504 42901 33507
rect 42852 33476 42901 33504
rect 42852 33464 42858 33476
rect 42889 33473 42901 33476
rect 42935 33473 42947 33507
rect 42889 33467 42947 33473
rect 42978 33464 42984 33516
rect 43036 33504 43042 33516
rect 43036 33476 43081 33504
rect 43036 33464 43042 33476
rect 46750 33464 46756 33516
rect 46808 33504 46814 33516
rect 46845 33507 46903 33513
rect 46845 33504 46857 33507
rect 46808 33476 46857 33504
rect 46808 33464 46814 33476
rect 46845 33473 46857 33476
rect 46891 33473 46903 33507
rect 46845 33467 46903 33473
rect 43622 33436 43628 33448
rect 40328 33408 40448 33436
rect 43583 33408 43628 33436
rect 40328 33380 40356 33408
rect 43622 33396 43628 33408
rect 43680 33396 43686 33448
rect 40310 33328 40316 33380
rect 40368 33328 40374 33380
rect 41230 33300 41236 33312
rect 40236 33272 41236 33300
rect 41230 33260 41236 33272
rect 41288 33260 41294 33312
rect 46934 33300 46940 33312
rect 46895 33272 46940 33300
rect 46934 33260 46940 33272
rect 46992 33260 46998 33312
rect 66254 33260 66260 33312
rect 66312 33300 66318 33312
rect 67637 33303 67695 33309
rect 67637 33300 67649 33303
rect 66312 33272 67649 33300
rect 66312 33260 66318 33272
rect 67637 33269 67649 33272
rect 67683 33269 67695 33303
rect 67637 33263 67695 33269
rect 1104 33210 68816 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 68816 33210
rect 1104 33136 68816 33158
rect 24946 33096 24952 33108
rect 24907 33068 24952 33096
rect 24946 33056 24952 33068
rect 25004 33056 25010 33108
rect 27614 33096 27620 33108
rect 27575 33068 27620 33096
rect 27614 33056 27620 33068
rect 27672 33056 27678 33108
rect 28166 33056 28172 33108
rect 28224 33096 28230 33108
rect 28261 33099 28319 33105
rect 28261 33096 28273 33099
rect 28224 33068 28273 33096
rect 28224 33056 28230 33068
rect 28261 33065 28273 33068
rect 28307 33065 28319 33099
rect 33778 33096 33784 33108
rect 33739 33068 33784 33096
rect 28261 33059 28319 33065
rect 33778 33056 33784 33068
rect 33836 33056 33842 33108
rect 34885 33099 34943 33105
rect 34885 33065 34897 33099
rect 34931 33096 34943 33099
rect 35710 33096 35716 33108
rect 34931 33068 35716 33096
rect 34931 33065 34943 33068
rect 34885 33059 34943 33065
rect 35710 33056 35716 33068
rect 35768 33056 35774 33108
rect 42886 33056 42892 33108
rect 42944 33096 42950 33108
rect 42981 33099 43039 33105
rect 42981 33096 42993 33099
rect 42944 33068 42993 33096
rect 42944 33056 42950 33068
rect 42981 33065 42993 33068
rect 43027 33065 43039 33099
rect 43622 33096 43628 33108
rect 43583 33068 43628 33096
rect 42981 33059 43039 33065
rect 43622 33056 43628 33068
rect 43680 33056 43686 33108
rect 36909 33031 36967 33037
rect 36909 32997 36921 33031
rect 36955 32997 36967 33031
rect 36909 32991 36967 32997
rect 23017 32895 23075 32901
rect 23017 32861 23029 32895
rect 23063 32892 23075 32895
rect 23382 32892 23388 32904
rect 23063 32864 23388 32892
rect 23063 32861 23075 32864
rect 23017 32855 23075 32861
rect 23382 32852 23388 32864
rect 23440 32852 23446 32904
rect 26234 32892 26240 32904
rect 26195 32864 26240 32892
rect 26234 32852 26240 32864
rect 26292 32852 26298 32904
rect 29638 32892 29644 32904
rect 26436 32864 29644 32892
rect 24857 32827 24915 32833
rect 24857 32793 24869 32827
rect 24903 32824 24915 32827
rect 25866 32824 25872 32836
rect 24903 32796 25872 32824
rect 24903 32793 24915 32796
rect 24857 32787 24915 32793
rect 25866 32784 25872 32796
rect 25924 32824 25930 32836
rect 26436 32824 26464 32864
rect 29638 32852 29644 32864
rect 29696 32852 29702 32904
rect 29733 32895 29791 32901
rect 29733 32861 29745 32895
rect 29779 32892 29791 32895
rect 29914 32892 29920 32904
rect 29779 32864 29920 32892
rect 29779 32861 29791 32864
rect 29733 32855 29791 32861
rect 29914 32852 29920 32864
rect 29972 32852 29978 32904
rect 31113 32895 31171 32901
rect 31113 32861 31125 32895
rect 31159 32892 31171 32895
rect 31386 32892 31392 32904
rect 31159 32864 31392 32892
rect 31159 32861 31171 32864
rect 31113 32855 31171 32861
rect 31386 32852 31392 32864
rect 31444 32852 31450 32904
rect 32398 32892 32404 32904
rect 32359 32864 32404 32892
rect 32398 32852 32404 32864
rect 32456 32852 32462 32904
rect 35529 32895 35587 32901
rect 35529 32861 35541 32895
rect 35575 32892 35587 32895
rect 35618 32892 35624 32904
rect 35575 32864 35624 32892
rect 35575 32861 35587 32864
rect 35529 32855 35587 32861
rect 35618 32852 35624 32864
rect 35676 32852 35682 32904
rect 36924 32892 36952 32991
rect 36998 32988 37004 33040
rect 37056 33028 37062 33040
rect 67266 33028 67272 33040
rect 37056 33000 67272 33028
rect 37056 32988 37062 33000
rect 67266 32988 67272 33000
rect 67324 32988 67330 33040
rect 37274 32920 37280 32972
rect 37332 32960 37338 32972
rect 46934 32960 46940 32972
rect 37332 32932 38700 32960
rect 46895 32932 46940 32960
rect 37332 32920 37338 32932
rect 37366 32892 37372 32904
rect 35728 32864 36952 32892
rect 37327 32864 37372 32892
rect 25924 32796 26464 32824
rect 26504 32827 26562 32833
rect 25924 32784 25930 32796
rect 26504 32793 26516 32827
rect 26550 32824 26562 32827
rect 26970 32824 26976 32836
rect 26550 32796 26976 32824
rect 26550 32793 26562 32796
rect 26504 32787 26562 32793
rect 26970 32784 26976 32796
rect 27028 32784 27034 32836
rect 27614 32784 27620 32836
rect 27672 32824 27678 32836
rect 28077 32827 28135 32833
rect 28077 32824 28089 32827
rect 27672 32796 28089 32824
rect 27672 32784 27678 32796
rect 28077 32793 28089 32796
rect 28123 32793 28135 32827
rect 28293 32827 28351 32833
rect 28293 32824 28305 32827
rect 28077 32787 28135 32793
rect 28184 32796 28305 32824
rect 22830 32756 22836 32768
rect 22791 32728 22836 32756
rect 22830 32716 22836 32728
rect 22888 32716 22894 32768
rect 27706 32716 27712 32768
rect 27764 32756 27770 32768
rect 28184 32756 28212 32796
rect 28293 32793 28305 32796
rect 28339 32824 28351 32827
rect 28810 32824 28816 32836
rect 28339 32796 28816 32824
rect 28339 32793 28351 32796
rect 28293 32787 28351 32793
rect 28810 32784 28816 32796
rect 28868 32784 28874 32836
rect 32668 32827 32726 32833
rect 32668 32793 32680 32827
rect 32714 32824 32726 32827
rect 32858 32824 32864 32836
rect 32714 32796 32864 32824
rect 32714 32793 32726 32796
rect 32668 32787 32726 32793
rect 32858 32784 32864 32796
rect 32916 32784 32922 32836
rect 33594 32784 33600 32836
rect 33652 32824 33658 32836
rect 34701 32827 34759 32833
rect 34701 32824 34713 32827
rect 33652 32796 34713 32824
rect 33652 32784 33658 32796
rect 34701 32793 34713 32796
rect 34747 32824 34759 32827
rect 35728 32824 35756 32864
rect 37366 32852 37372 32864
rect 37424 32852 37430 32904
rect 37458 32852 37464 32904
rect 37516 32892 37522 32904
rect 38672 32901 38700 32932
rect 46934 32920 46940 32932
rect 46992 32920 46998 32972
rect 66254 32960 66260 32972
rect 66215 32932 66260 32960
rect 66254 32920 66260 32932
rect 66312 32920 66318 32972
rect 37553 32895 37611 32901
rect 37553 32892 37565 32895
rect 37516 32864 37565 32892
rect 37516 32852 37522 32864
rect 37553 32861 37565 32864
rect 37599 32861 37611 32895
rect 37553 32855 37611 32861
rect 38657 32895 38715 32901
rect 38657 32861 38669 32895
rect 38703 32861 38715 32895
rect 38657 32855 38715 32861
rect 42426 32852 42432 32904
rect 42484 32892 42490 32904
rect 42613 32895 42671 32901
rect 42613 32892 42625 32895
rect 42484 32864 42625 32892
rect 42484 32852 42490 32864
rect 42613 32861 42625 32864
rect 42659 32861 42671 32895
rect 42794 32892 42800 32904
rect 42755 32864 42800 32892
rect 42613 32855 42671 32861
rect 42794 32852 42800 32864
rect 42852 32852 42858 32904
rect 43438 32892 43444 32904
rect 43399 32864 43444 32892
rect 43438 32852 43444 32864
rect 43496 32852 43502 32904
rect 44266 32892 44272 32904
rect 44227 32864 44272 32892
rect 44266 32852 44272 32864
rect 44324 32852 44330 32904
rect 46750 32892 46756 32904
rect 46711 32864 46756 32892
rect 46750 32852 46756 32864
rect 46808 32852 46814 32904
rect 34747 32796 35756 32824
rect 35796 32827 35854 32833
rect 34747 32793 34759 32796
rect 34701 32787 34759 32793
rect 35796 32793 35808 32827
rect 35842 32824 35854 32827
rect 36446 32824 36452 32836
rect 35842 32796 36452 32824
rect 35842 32793 35854 32796
rect 35796 32787 35854 32793
rect 36446 32784 36452 32796
rect 36504 32784 36510 32836
rect 48593 32827 48651 32833
rect 48593 32793 48605 32827
rect 48639 32824 48651 32827
rect 65518 32824 65524 32836
rect 48639 32796 65524 32824
rect 48639 32793 48651 32796
rect 48593 32787 48651 32793
rect 65518 32784 65524 32796
rect 65576 32784 65582 32836
rect 66438 32824 66444 32836
rect 66399 32796 66444 32824
rect 66438 32784 66444 32796
rect 66496 32784 66502 32836
rect 68094 32824 68100 32836
rect 68055 32796 68100 32824
rect 68094 32784 68100 32796
rect 68152 32784 68158 32836
rect 28442 32756 28448 32768
rect 27764 32728 28212 32756
rect 28403 32728 28448 32756
rect 27764 32716 27770 32728
rect 28442 32716 28448 32728
rect 28500 32716 28506 32768
rect 29546 32756 29552 32768
rect 29507 32728 29552 32756
rect 29546 32716 29552 32728
rect 29604 32716 29610 32768
rect 30834 32716 30840 32768
rect 30892 32756 30898 32768
rect 30929 32759 30987 32765
rect 30929 32756 30941 32759
rect 30892 32728 30941 32756
rect 30892 32716 30898 32728
rect 30929 32725 30941 32728
rect 30975 32725 30987 32759
rect 30929 32719 30987 32725
rect 34882 32716 34888 32768
rect 34940 32765 34946 32768
rect 34940 32759 34959 32765
rect 34947 32725 34959 32759
rect 34940 32719 34959 32725
rect 35069 32759 35127 32765
rect 35069 32725 35081 32759
rect 35115 32756 35127 32759
rect 36630 32756 36636 32768
rect 35115 32728 36636 32756
rect 35115 32725 35127 32728
rect 35069 32719 35127 32725
rect 34940 32716 34946 32719
rect 36630 32716 36636 32728
rect 36688 32716 36694 32768
rect 37737 32759 37795 32765
rect 37737 32725 37749 32759
rect 37783 32756 37795 32759
rect 38378 32756 38384 32768
rect 37783 32728 38384 32756
rect 37783 32725 37795 32728
rect 37737 32719 37795 32725
rect 38378 32716 38384 32728
rect 38436 32716 38442 32768
rect 38749 32759 38807 32765
rect 38749 32725 38761 32759
rect 38795 32756 38807 32759
rect 39298 32756 39304 32768
rect 38795 32728 39304 32756
rect 38795 32725 38807 32728
rect 38749 32719 38807 32725
rect 39298 32716 39304 32728
rect 39356 32716 39362 32768
rect 43714 32716 43720 32768
rect 43772 32756 43778 32768
rect 44361 32759 44419 32765
rect 44361 32756 44373 32759
rect 43772 32728 44373 32756
rect 43772 32716 43778 32728
rect 44361 32725 44373 32728
rect 44407 32725 44419 32759
rect 44361 32719 44419 32725
rect 1104 32666 68816 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 68816 32666
rect 1104 32592 68816 32614
rect 25314 32512 25320 32564
rect 25372 32552 25378 32564
rect 25685 32555 25743 32561
rect 25685 32552 25697 32555
rect 25372 32524 25697 32552
rect 25372 32512 25378 32524
rect 25685 32521 25697 32524
rect 25731 32521 25743 32555
rect 25685 32515 25743 32521
rect 26234 32512 26240 32564
rect 26292 32552 26298 32564
rect 26329 32555 26387 32561
rect 26329 32552 26341 32555
rect 26292 32524 26341 32552
rect 26292 32512 26298 32524
rect 26329 32521 26341 32524
rect 26375 32521 26387 32555
rect 26970 32552 26976 32564
rect 26931 32524 26976 32552
rect 26329 32515 26387 32521
rect 26970 32512 26976 32524
rect 27028 32512 27034 32564
rect 29638 32512 29644 32564
rect 29696 32552 29702 32564
rect 30098 32552 30104 32564
rect 29696 32524 30104 32552
rect 29696 32512 29702 32524
rect 30098 32512 30104 32524
rect 30156 32512 30162 32564
rect 31386 32552 31392 32564
rect 31347 32524 31392 32552
rect 31386 32512 31392 32524
rect 31444 32512 31450 32564
rect 32398 32552 32404 32564
rect 32359 32524 32404 32552
rect 32398 32512 32404 32524
rect 32456 32512 32462 32564
rect 34882 32512 34888 32564
rect 34940 32552 34946 32564
rect 35802 32552 35808 32564
rect 34940 32524 35808 32552
rect 34940 32512 34946 32524
rect 35802 32512 35808 32524
rect 35860 32512 35866 32564
rect 36446 32552 36452 32564
rect 36407 32524 36452 32552
rect 36446 32512 36452 32524
rect 36504 32512 36510 32564
rect 44085 32555 44143 32561
rect 44085 32521 44097 32555
rect 44131 32552 44143 32555
rect 44131 32524 45692 32552
rect 44131 32521 44143 32524
rect 44085 32515 44143 32521
rect 22640 32487 22698 32493
rect 22640 32453 22652 32487
rect 22686 32484 22698 32487
rect 22830 32484 22836 32496
rect 22686 32456 22836 32484
rect 22686 32453 22698 32456
rect 22640 32447 22698 32453
rect 22830 32444 22836 32456
rect 22888 32444 22894 32496
rect 25774 32484 25780 32496
rect 25424 32456 25780 32484
rect 25424 32425 25452 32456
rect 25774 32444 25780 32456
rect 25832 32444 25838 32496
rect 28988 32487 29046 32493
rect 28988 32453 29000 32487
rect 29034 32484 29046 32487
rect 29546 32484 29552 32496
rect 29034 32456 29552 32484
rect 29034 32453 29046 32456
rect 28988 32447 29046 32453
rect 29546 32444 29552 32456
rect 29604 32444 29610 32496
rect 35253 32487 35311 32493
rect 35253 32453 35265 32487
rect 35299 32484 35311 32487
rect 37277 32487 37335 32493
rect 37277 32484 37289 32487
rect 35299 32456 37289 32484
rect 35299 32453 35311 32456
rect 35253 32447 35311 32453
rect 37277 32453 37289 32456
rect 37323 32453 37335 32487
rect 37277 32447 37335 32453
rect 37366 32444 37372 32496
rect 37424 32484 37430 32496
rect 37461 32487 37519 32493
rect 37461 32484 37473 32487
rect 37424 32456 37473 32484
rect 37424 32444 37430 32456
rect 37461 32453 37473 32456
rect 37507 32484 37519 32487
rect 37642 32484 37648 32496
rect 37507 32456 37648 32484
rect 37507 32453 37519 32456
rect 37461 32447 37519 32453
rect 37642 32444 37648 32456
rect 37700 32444 37706 32496
rect 39390 32484 39396 32496
rect 38580 32456 39396 32484
rect 25409 32419 25467 32425
rect 25409 32385 25421 32419
rect 25455 32385 25467 32419
rect 25409 32379 25467 32385
rect 25498 32376 25504 32428
rect 25556 32416 25562 32428
rect 25556 32388 25601 32416
rect 25556 32376 25562 32388
rect 26050 32376 26056 32428
rect 26108 32416 26114 32428
rect 26145 32419 26203 32425
rect 26145 32416 26157 32419
rect 26108 32388 26157 32416
rect 26108 32376 26114 32388
rect 26145 32385 26157 32388
rect 26191 32385 26203 32419
rect 26145 32379 26203 32385
rect 27157 32419 27215 32425
rect 27157 32385 27169 32419
rect 27203 32416 27215 32419
rect 28442 32416 28448 32428
rect 27203 32388 28448 32416
rect 27203 32385 27215 32388
rect 27157 32379 27215 32385
rect 28442 32376 28448 32388
rect 28500 32376 28506 32428
rect 31205 32419 31263 32425
rect 31205 32385 31217 32419
rect 31251 32416 31263 32419
rect 31294 32416 31300 32428
rect 31251 32388 31300 32416
rect 31251 32385 31263 32388
rect 31205 32379 31263 32385
rect 31294 32376 31300 32388
rect 31352 32416 31358 32428
rect 31846 32416 31852 32428
rect 31352 32388 31852 32416
rect 31352 32376 31358 32388
rect 31846 32376 31852 32388
rect 31904 32376 31910 32428
rect 32306 32416 32312 32428
rect 32267 32388 32312 32416
rect 32306 32376 32312 32388
rect 32364 32376 32370 32428
rect 33413 32419 33471 32425
rect 33413 32385 33425 32419
rect 33459 32416 33471 32419
rect 33778 32416 33784 32428
rect 33459 32388 33784 32416
rect 33459 32385 33471 32388
rect 33413 32379 33471 32385
rect 33778 32376 33784 32388
rect 33836 32376 33842 32428
rect 35434 32376 35440 32428
rect 35492 32416 35498 32428
rect 35805 32419 35863 32425
rect 35805 32416 35817 32419
rect 35492 32388 35817 32416
rect 35492 32376 35498 32388
rect 35805 32385 35817 32388
rect 35851 32385 35863 32419
rect 36630 32416 36636 32428
rect 36591 32388 36636 32416
rect 35805 32379 35863 32385
rect 36630 32376 36636 32388
rect 36688 32376 36694 32428
rect 38378 32416 38384 32428
rect 38339 32388 38384 32416
rect 38378 32376 38384 32388
rect 38436 32376 38442 32428
rect 38580 32425 38608 32456
rect 39390 32444 39396 32456
rect 39448 32444 39454 32496
rect 39482 32444 39488 32496
rect 39540 32444 39546 32496
rect 42610 32444 42616 32496
rect 42668 32484 42674 32496
rect 42889 32487 42947 32493
rect 42889 32484 42901 32487
rect 42668 32456 42901 32484
rect 42668 32444 42674 32456
rect 42889 32453 42901 32456
rect 42935 32453 42947 32487
rect 42889 32447 42947 32453
rect 43714 32444 43720 32496
rect 43772 32484 43778 32496
rect 45554 32484 45560 32496
rect 43772 32456 44772 32484
rect 43772 32444 43778 32456
rect 38565 32419 38623 32425
rect 38565 32385 38577 32419
rect 38611 32385 38623 32419
rect 39298 32416 39304 32428
rect 39259 32388 39304 32416
rect 38565 32379 38623 32385
rect 39298 32376 39304 32388
rect 39356 32376 39362 32428
rect 39500 32416 39528 32444
rect 39574 32425 39580 32428
rect 39408 32388 39528 32416
rect 22370 32348 22376 32360
rect 22331 32320 22376 32348
rect 22370 32308 22376 32320
rect 22428 32308 22434 32360
rect 28718 32348 28724 32360
rect 28679 32320 28724 32348
rect 28718 32308 28724 32320
rect 28776 32308 28782 32360
rect 31021 32351 31079 32357
rect 31021 32317 31033 32351
rect 31067 32348 31079 32351
rect 31938 32348 31944 32360
rect 31067 32320 31944 32348
rect 31067 32317 31079 32320
rect 31021 32311 31079 32317
rect 31938 32308 31944 32320
rect 31996 32308 32002 32360
rect 33594 32348 33600 32360
rect 33555 32320 33600 32348
rect 33594 32308 33600 32320
rect 33652 32308 33658 32360
rect 34333 32351 34391 32357
rect 34333 32348 34345 32351
rect 33704 32320 34345 32348
rect 23753 32283 23811 32289
rect 23753 32249 23765 32283
rect 23799 32280 23811 32283
rect 28258 32280 28264 32292
rect 23799 32252 28264 32280
rect 23799 32249 23811 32252
rect 23753 32243 23811 32249
rect 23014 32172 23020 32224
rect 23072 32212 23078 32224
rect 23768 32212 23796 32243
rect 28258 32240 28264 32252
rect 28316 32240 28322 32292
rect 32950 32240 32956 32292
rect 33008 32280 33014 32292
rect 33704 32280 33732 32320
rect 34333 32317 34345 32320
rect 34379 32317 34391 32351
rect 34333 32311 34391 32317
rect 34422 32308 34428 32360
rect 34480 32357 34486 32360
rect 34480 32351 34508 32357
rect 34496 32317 34508 32351
rect 34480 32311 34508 32317
rect 34609 32351 34667 32357
rect 34609 32317 34621 32351
rect 34655 32348 34667 32351
rect 35342 32348 35348 32360
rect 34655 32320 35348 32348
rect 34655 32317 34667 32320
rect 34609 32311 34667 32317
rect 34480 32308 34486 32311
rect 35342 32308 35348 32320
rect 35400 32308 35406 32360
rect 38286 32348 38292 32360
rect 38247 32320 38292 32348
rect 38286 32308 38292 32320
rect 38344 32308 38350 32360
rect 38473 32351 38531 32357
rect 38473 32317 38485 32351
rect 38519 32348 38531 32351
rect 39408 32348 39436 32388
rect 39568 32379 39580 32425
rect 39632 32416 39638 32428
rect 39632 32388 39668 32416
rect 39574 32376 39580 32379
rect 39632 32376 39638 32388
rect 41138 32376 41144 32428
rect 41196 32416 41202 32428
rect 41233 32419 41291 32425
rect 41233 32416 41245 32419
rect 41196 32388 41245 32416
rect 41196 32376 41202 32388
rect 41233 32385 41245 32388
rect 41279 32385 41291 32419
rect 41233 32379 41291 32385
rect 42426 32376 42432 32428
rect 42484 32416 42490 32428
rect 42702 32416 42708 32428
rect 42484 32388 42708 32416
rect 42484 32376 42490 32388
rect 42702 32376 42708 32388
rect 42760 32376 42766 32428
rect 43070 32376 43076 32428
rect 43128 32416 43134 32428
rect 43622 32416 43628 32428
rect 43128 32388 43628 32416
rect 43128 32376 43134 32388
rect 43622 32376 43628 32388
rect 43680 32376 43686 32428
rect 44358 32416 44364 32428
rect 44319 32388 44364 32416
rect 44358 32376 44364 32388
rect 44416 32376 44422 32428
rect 44450 32419 44508 32425
rect 44450 32385 44462 32419
rect 44496 32385 44508 32419
rect 44450 32379 44508 32385
rect 38519 32320 39436 32348
rect 38519 32317 38531 32320
rect 38473 32311 38531 32317
rect 41322 32308 41328 32360
rect 41380 32348 41386 32360
rect 44468 32348 44496 32379
rect 44542 32376 44548 32428
rect 44600 32416 44606 32428
rect 44744 32425 44772 32456
rect 45204 32456 45560 32484
rect 44729 32419 44787 32425
rect 44600 32388 44645 32416
rect 44600 32376 44606 32388
rect 44729 32385 44741 32419
rect 44775 32385 44787 32419
rect 44729 32379 44787 32385
rect 44634 32348 44640 32360
rect 41380 32320 44312 32348
rect 44468 32320 44640 32348
rect 41380 32308 41386 32320
rect 34054 32280 34060 32292
rect 33008 32252 33732 32280
rect 34015 32252 34060 32280
rect 33008 32240 33014 32252
rect 34054 32240 34060 32252
rect 34112 32240 34118 32292
rect 37645 32283 37703 32289
rect 37645 32249 37657 32283
rect 37691 32280 37703 32283
rect 42058 32280 42064 32292
rect 37691 32252 39344 32280
rect 37691 32249 37703 32252
rect 37645 32243 37703 32249
rect 35894 32212 35900 32224
rect 23072 32184 23796 32212
rect 35855 32184 35900 32212
rect 23072 32172 23078 32184
rect 35894 32172 35900 32184
rect 35952 32172 35958 32224
rect 38102 32212 38108 32224
rect 38063 32184 38108 32212
rect 38102 32172 38108 32184
rect 38160 32172 38166 32224
rect 39316 32212 39344 32252
rect 40236 32252 42064 32280
rect 40236 32212 40264 32252
rect 42058 32240 42064 32252
rect 42116 32240 42122 32292
rect 44284 32280 44312 32320
rect 44634 32308 44640 32320
rect 44692 32308 44698 32360
rect 45204 32357 45232 32456
rect 45554 32444 45560 32456
rect 45612 32444 45618 32496
rect 45456 32419 45514 32425
rect 45456 32385 45468 32419
rect 45502 32416 45514 32419
rect 45664 32416 45692 32524
rect 66438 32512 66444 32564
rect 66496 32552 66502 32564
rect 67545 32555 67603 32561
rect 67545 32552 67557 32555
rect 66496 32524 67557 32552
rect 66496 32512 66502 32524
rect 67545 32521 67557 32524
rect 67591 32521 67603 32555
rect 67545 32515 67603 32521
rect 45502 32388 45692 32416
rect 45502 32385 45514 32388
rect 45456 32379 45514 32385
rect 67266 32376 67272 32428
rect 67324 32416 67330 32428
rect 67453 32419 67511 32425
rect 67453 32416 67465 32419
rect 67324 32388 67465 32416
rect 67324 32376 67330 32388
rect 67453 32385 67465 32388
rect 67499 32385 67511 32419
rect 67453 32379 67511 32385
rect 45189 32351 45247 32357
rect 45189 32317 45201 32351
rect 45235 32317 45247 32351
rect 45189 32311 45247 32317
rect 45204 32280 45232 32311
rect 44284 32252 45232 32280
rect 40678 32212 40684 32224
rect 39316 32184 40264 32212
rect 40639 32184 40684 32212
rect 40678 32172 40684 32184
rect 40736 32172 40742 32224
rect 41322 32172 41328 32224
rect 41380 32212 41386 32224
rect 41417 32215 41475 32221
rect 41417 32212 41429 32215
rect 41380 32184 41429 32212
rect 41380 32172 41386 32184
rect 41417 32181 41429 32184
rect 41463 32181 41475 32215
rect 41417 32175 41475 32181
rect 43073 32215 43131 32221
rect 43073 32181 43085 32215
rect 43119 32212 43131 32215
rect 43346 32212 43352 32224
rect 43119 32184 43352 32212
rect 43119 32181 43131 32184
rect 43073 32175 43131 32181
rect 43346 32172 43352 32184
rect 43404 32172 43410 32224
rect 44358 32172 44364 32224
rect 44416 32212 44422 32224
rect 46569 32215 46627 32221
rect 46569 32212 46581 32215
rect 44416 32184 46581 32212
rect 44416 32172 44422 32184
rect 46569 32181 46581 32184
rect 46615 32212 46627 32215
rect 46750 32212 46756 32224
rect 46615 32184 46756 32212
rect 46615 32181 46627 32184
rect 46569 32175 46627 32181
rect 46750 32172 46756 32184
rect 46808 32172 46814 32224
rect 1104 32122 68816 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 68816 32122
rect 1104 32048 68816 32070
rect 22370 31968 22376 32020
rect 22428 32008 22434 32020
rect 22465 32011 22523 32017
rect 22465 32008 22477 32011
rect 22428 31980 22477 32008
rect 22428 31968 22434 31980
rect 22465 31977 22477 31980
rect 22511 31977 22523 32011
rect 23382 32008 23388 32020
rect 23343 31980 23388 32008
rect 22465 31971 22523 31977
rect 23382 31968 23388 31980
rect 23440 31968 23446 32020
rect 28718 31968 28724 32020
rect 28776 32008 28782 32020
rect 28813 32011 28871 32017
rect 28813 32008 28825 32011
rect 28776 31980 28825 32008
rect 28776 31968 28782 31980
rect 28813 31977 28825 31980
rect 28859 31977 28871 32011
rect 28813 31971 28871 31977
rect 29086 31968 29092 32020
rect 29144 32008 29150 32020
rect 29733 32011 29791 32017
rect 29733 32008 29745 32011
rect 29144 31980 29745 32008
rect 29144 31968 29150 31980
rect 29733 31977 29745 31980
rect 29779 31977 29791 32011
rect 29914 32008 29920 32020
rect 29875 31980 29920 32008
rect 29733 31971 29791 31977
rect 29914 31968 29920 31980
rect 29972 31968 29978 32020
rect 32858 32008 32864 32020
rect 32819 31980 32864 32008
rect 32858 31968 32864 31980
rect 32916 31968 32922 32020
rect 35618 32008 35624 32020
rect 35579 31980 35624 32008
rect 35618 31968 35624 31980
rect 35676 31968 35682 32020
rect 38286 31968 38292 32020
rect 38344 32008 38350 32020
rect 39209 32011 39267 32017
rect 39209 32008 39221 32011
rect 38344 31980 39221 32008
rect 38344 31968 38350 31980
rect 39209 31977 39221 31980
rect 39255 31977 39267 32011
rect 39209 31971 39267 31977
rect 43165 32011 43223 32017
rect 43165 31977 43177 32011
rect 43211 32008 43223 32011
rect 44542 32008 44548 32020
rect 43211 31980 44548 32008
rect 43211 31977 43223 31980
rect 43165 31971 43223 31977
rect 44542 31968 44548 31980
rect 44600 31968 44606 32020
rect 31938 31940 31944 31952
rect 31851 31912 31944 31940
rect 31938 31900 31944 31912
rect 31996 31940 32002 31952
rect 34422 31940 34428 31952
rect 31996 31912 34428 31940
rect 31996 31900 32002 31912
rect 34422 31900 34428 31912
rect 34480 31900 34486 31952
rect 37277 31943 37335 31949
rect 37277 31909 37289 31943
rect 37323 31940 37335 31943
rect 37323 31912 40816 31940
rect 37323 31909 37335 31912
rect 37277 31903 37335 31909
rect 23014 31872 23020 31884
rect 22975 31844 23020 31872
rect 23014 31832 23020 31844
rect 23072 31832 23078 31884
rect 23566 31872 23572 31884
rect 23216 31844 23572 31872
rect 1670 31764 1676 31816
rect 1728 31804 1734 31816
rect 1857 31807 1915 31813
rect 1857 31804 1869 31807
rect 1728 31776 1869 31804
rect 1728 31764 1734 31776
rect 1857 31773 1869 31776
rect 1903 31773 1915 31807
rect 22462 31804 22468 31816
rect 22423 31776 22468 31804
rect 1857 31767 1915 31773
rect 22462 31764 22468 31776
rect 22520 31764 22526 31816
rect 23216 31813 23244 31844
rect 23566 31832 23572 31844
rect 23624 31872 23630 31884
rect 24765 31875 24823 31881
rect 24765 31872 24777 31875
rect 23624 31844 24777 31872
rect 23624 31832 23630 31844
rect 24765 31841 24777 31844
rect 24811 31841 24823 31875
rect 27798 31872 27804 31884
rect 24765 31835 24823 31841
rect 25884 31844 27804 31872
rect 23201 31807 23259 31813
rect 23201 31773 23213 31807
rect 23247 31773 23259 31807
rect 23201 31767 23259 31773
rect 24489 31807 24547 31813
rect 24489 31773 24501 31807
rect 24535 31804 24547 31807
rect 25884 31804 25912 31844
rect 27798 31832 27804 31844
rect 27856 31872 27862 31884
rect 28902 31872 28908 31884
rect 27856 31844 28908 31872
rect 27856 31832 27862 31844
rect 28902 31832 28908 31844
rect 28960 31832 28966 31884
rect 29730 31832 29736 31884
rect 29788 31832 29794 31884
rect 30558 31872 30564 31884
rect 30519 31844 30564 31872
rect 30558 31832 30564 31844
rect 30616 31832 30622 31884
rect 33962 31832 33968 31884
rect 34020 31872 34026 31884
rect 39853 31875 39911 31881
rect 39853 31872 39865 31875
rect 34020 31844 36952 31872
rect 34020 31832 34026 31844
rect 24535 31776 25912 31804
rect 25961 31807 26019 31813
rect 24535 31773 24547 31776
rect 24489 31767 24547 31773
rect 25961 31773 25973 31807
rect 26007 31804 26019 31807
rect 26050 31804 26056 31816
rect 26007 31776 26056 31804
rect 26007 31773 26019 31776
rect 25961 31767 26019 31773
rect 26050 31764 26056 31776
rect 26108 31764 26114 31816
rect 26694 31804 26700 31816
rect 26655 31776 26700 31804
rect 26694 31764 26700 31776
rect 26752 31764 26758 31816
rect 28534 31764 28540 31816
rect 28592 31804 28598 31816
rect 28629 31807 28687 31813
rect 28629 31804 28641 31807
rect 28592 31776 28641 31804
rect 28592 31764 28598 31776
rect 28629 31773 28641 31776
rect 28675 31773 28687 31807
rect 28629 31767 28687 31773
rect 29764 31754 29792 31832
rect 30834 31813 30840 31816
rect 30828 31804 30840 31813
rect 30795 31776 30840 31804
rect 30828 31767 30840 31776
rect 30834 31764 30840 31767
rect 30892 31764 30898 31816
rect 33045 31807 33103 31813
rect 33045 31773 33057 31807
rect 33091 31804 33103 31807
rect 33318 31804 33324 31816
rect 33091 31776 33324 31804
rect 33091 31773 33103 31776
rect 33045 31767 33103 31773
rect 33318 31764 33324 31776
rect 33376 31764 33382 31816
rect 35621 31807 35679 31813
rect 35621 31773 35633 31807
rect 35667 31804 35679 31807
rect 35710 31804 35716 31816
rect 35667 31776 35716 31804
rect 35667 31773 35679 31776
rect 35621 31767 35679 31773
rect 35710 31764 35716 31776
rect 35768 31764 35774 31816
rect 36924 31813 36952 31844
rect 39040 31844 39865 31872
rect 36909 31807 36967 31813
rect 36909 31773 36921 31807
rect 36955 31773 36967 31807
rect 36909 31767 36967 31773
rect 37093 31807 37151 31813
rect 37093 31773 37105 31807
rect 37139 31804 37151 31807
rect 37366 31804 37372 31816
rect 37139 31776 37372 31804
rect 37139 31773 37151 31776
rect 37093 31767 37151 31773
rect 37366 31764 37372 31776
rect 37424 31764 37430 31816
rect 38838 31804 38844 31816
rect 38799 31776 38844 31804
rect 38838 31764 38844 31776
rect 38896 31764 38902 31816
rect 39040 31813 39068 31844
rect 39853 31841 39865 31844
rect 39899 31872 39911 31875
rect 40678 31872 40684 31884
rect 39899 31844 40684 31872
rect 39899 31841 39911 31844
rect 39853 31835 39911 31841
rect 40678 31832 40684 31844
rect 40736 31832 40742 31884
rect 39025 31807 39083 31813
rect 39025 31773 39037 31807
rect 39071 31773 39083 31807
rect 40034 31804 40040 31816
rect 39995 31776 40040 31804
rect 39025 31767 39083 31773
rect 40034 31764 40040 31776
rect 40092 31764 40098 31816
rect 40788 31804 40816 31912
rect 42610 31900 42616 31952
rect 42668 31940 42674 31952
rect 42705 31943 42763 31949
rect 42705 31940 42717 31943
rect 42668 31912 42717 31940
rect 42668 31900 42674 31912
rect 42705 31909 42717 31912
rect 42751 31909 42763 31943
rect 42705 31903 42763 31909
rect 43254 31900 43260 31952
rect 43312 31940 43318 31952
rect 43312 31912 43576 31940
rect 43312 31900 43318 31912
rect 41322 31872 41328 31884
rect 41283 31844 41328 31872
rect 41322 31832 41328 31844
rect 41380 31832 41386 31884
rect 43548 31881 43576 31912
rect 43441 31875 43499 31881
rect 43441 31872 43453 31875
rect 43272 31844 43453 31872
rect 43272 31804 43300 31844
rect 43441 31841 43453 31844
rect 43487 31841 43499 31875
rect 43441 31835 43499 31841
rect 43533 31875 43591 31881
rect 43533 31841 43545 31875
rect 43579 31841 43591 31875
rect 43533 31835 43591 31841
rect 43622 31832 43628 31884
rect 43680 31872 43686 31884
rect 43680 31844 43725 31872
rect 43680 31832 43686 31844
rect 40788 31776 43300 31804
rect 43346 31764 43352 31816
rect 43404 31804 43410 31816
rect 43404 31776 43449 31804
rect 43404 31764 43410 31776
rect 66254 31764 66260 31816
rect 66312 31804 66318 31816
rect 67913 31807 67971 31813
rect 67913 31804 67925 31807
rect 66312 31776 67925 31804
rect 66312 31764 66318 31776
rect 67913 31773 67925 31776
rect 67959 31773 67971 31807
rect 67913 31767 67971 31773
rect 29748 31748 29792 31754
rect 29549 31739 29607 31745
rect 29549 31705 29561 31739
rect 29595 31736 29607 31739
rect 29638 31736 29644 31748
rect 29595 31708 29644 31736
rect 29595 31705 29607 31708
rect 29549 31699 29607 31705
rect 29638 31696 29644 31708
rect 29696 31696 29702 31748
rect 29730 31696 29736 31748
rect 29788 31745 29794 31748
rect 29788 31739 29807 31745
rect 29795 31736 29807 31739
rect 29795 31708 29881 31736
rect 29795 31705 29807 31708
rect 29788 31699 29807 31705
rect 29788 31696 29794 31699
rect 37826 31696 37832 31748
rect 37884 31736 37890 31748
rect 41138 31736 41144 31748
rect 37884 31708 41144 31736
rect 37884 31696 37890 31708
rect 41138 31696 41144 31708
rect 41196 31696 41202 31748
rect 41592 31739 41650 31745
rect 41592 31705 41604 31739
rect 41638 31736 41650 31739
rect 41690 31736 41696 31748
rect 41638 31708 41696 31736
rect 41638 31705 41650 31708
rect 41592 31699 41650 31705
rect 41690 31696 41696 31708
rect 41748 31696 41754 31748
rect 25038 31628 25044 31680
rect 25096 31668 25102 31680
rect 25961 31671 26019 31677
rect 25961 31668 25973 31671
rect 25096 31640 25973 31668
rect 25096 31628 25102 31640
rect 25961 31637 25973 31640
rect 26007 31637 26019 31671
rect 26510 31668 26516 31680
rect 26471 31640 26516 31668
rect 25961 31631 26019 31637
rect 26510 31628 26516 31640
rect 26568 31628 26574 31680
rect 34698 31628 34704 31680
rect 34756 31668 34762 31680
rect 35618 31668 35624 31680
rect 34756 31640 35624 31668
rect 34756 31628 34762 31640
rect 35618 31628 35624 31640
rect 35676 31628 35682 31680
rect 40218 31668 40224 31680
rect 40179 31640 40224 31668
rect 40218 31628 40224 31640
rect 40276 31628 40282 31680
rect 41156 31668 41184 31696
rect 43438 31668 43444 31680
rect 41156 31640 43444 31668
rect 43438 31628 43444 31640
rect 43496 31628 43502 31680
rect 1104 31578 68816 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 68816 31578
rect 1104 31504 68816 31526
rect 22462 31424 22468 31476
rect 22520 31464 22526 31476
rect 23198 31464 23204 31476
rect 22520 31436 23204 31464
rect 22520 31424 22526 31436
rect 23198 31424 23204 31436
rect 23256 31424 23262 31476
rect 26694 31424 26700 31476
rect 26752 31464 26758 31476
rect 27341 31467 27399 31473
rect 27341 31464 27353 31467
rect 26752 31436 27353 31464
rect 26752 31424 26758 31436
rect 27341 31433 27353 31436
rect 27387 31433 27399 31467
rect 27341 31427 27399 31433
rect 27706 31424 27712 31476
rect 27764 31464 27770 31476
rect 28001 31467 28059 31473
rect 28001 31464 28013 31467
rect 27764 31436 28013 31464
rect 27764 31424 27770 31436
rect 28001 31433 28013 31436
rect 28047 31433 28059 31467
rect 28001 31427 28059 31433
rect 39574 31424 39580 31476
rect 39632 31464 39638 31476
rect 39669 31467 39727 31473
rect 39669 31464 39681 31467
rect 39632 31436 39681 31464
rect 39632 31424 39638 31436
rect 39669 31433 39681 31436
rect 39715 31433 39727 31467
rect 41690 31464 41696 31476
rect 41651 31436 41696 31464
rect 39669 31427 39727 31433
rect 41690 31424 41696 31436
rect 41748 31424 41754 31476
rect 25308 31399 25366 31405
rect 25308 31365 25320 31399
rect 25354 31396 25366 31399
rect 26510 31396 26516 31408
rect 25354 31368 26516 31396
rect 25354 31365 25366 31368
rect 25308 31359 25366 31365
rect 26510 31356 26516 31368
rect 26568 31356 26574 31408
rect 26973 31399 27031 31405
rect 26973 31365 26985 31399
rect 27019 31365 27031 31399
rect 26973 31359 27031 31365
rect 27189 31399 27247 31405
rect 27189 31365 27201 31399
rect 27235 31396 27247 31399
rect 27724 31396 27752 31424
rect 27235 31368 27752 31396
rect 27235 31365 27247 31368
rect 27189 31359 27247 31365
rect 1670 31328 1676 31340
rect 1631 31300 1676 31328
rect 1670 31288 1676 31300
rect 1728 31288 1734 31340
rect 23017 31331 23075 31337
rect 23017 31297 23029 31331
rect 23063 31297 23075 31331
rect 25038 31328 25044 31340
rect 24999 31300 25044 31328
rect 23017 31291 23075 31297
rect 1857 31263 1915 31269
rect 1857 31229 1869 31263
rect 1903 31260 1915 31263
rect 2038 31260 2044 31272
rect 1903 31232 2044 31260
rect 1903 31229 1915 31232
rect 1857 31223 1915 31229
rect 2038 31220 2044 31232
rect 2096 31220 2102 31272
rect 2774 31260 2780 31272
rect 2735 31232 2780 31260
rect 2774 31220 2780 31232
rect 2832 31220 2838 31272
rect 23032 31192 23060 31291
rect 25038 31288 25044 31300
rect 25096 31288 25102 31340
rect 26988 31328 27016 31359
rect 27798 31356 27804 31408
rect 27856 31396 27862 31408
rect 27856 31368 27901 31396
rect 27856 31356 27862 31368
rect 34514 31356 34520 31408
rect 34572 31396 34578 31408
rect 35345 31399 35403 31405
rect 35345 31396 35357 31399
rect 34572 31368 35357 31396
rect 34572 31356 34578 31368
rect 35345 31365 35357 31368
rect 35391 31365 35403 31399
rect 35345 31359 35403 31365
rect 35434 31356 35440 31408
rect 35492 31396 35498 31408
rect 35545 31399 35603 31405
rect 35545 31396 35557 31399
rect 35492 31368 35557 31396
rect 35492 31356 35498 31368
rect 35545 31365 35557 31368
rect 35591 31396 35603 31399
rect 35802 31396 35808 31408
rect 35591 31368 35808 31396
rect 35591 31365 35603 31368
rect 35545 31359 35603 31365
rect 35802 31356 35808 31368
rect 35860 31356 35866 31408
rect 38838 31396 38844 31408
rect 38751 31368 38844 31396
rect 38838 31356 38844 31368
rect 38896 31396 38902 31408
rect 39206 31396 39212 31408
rect 38896 31368 39212 31396
rect 38896 31356 38902 31368
rect 39206 31356 39212 31368
rect 39264 31356 39270 31408
rect 66254 31396 66260 31408
rect 65812 31368 66260 31396
rect 26528 31300 27016 31328
rect 31573 31331 31631 31337
rect 23032 31164 24624 31192
rect 24596 31124 24624 31164
rect 26528 31136 26556 31300
rect 31573 31297 31585 31331
rect 31619 31328 31631 31331
rect 32214 31328 32220 31340
rect 31619 31300 32220 31328
rect 31619 31297 31631 31300
rect 31573 31291 31631 31297
rect 32214 31288 32220 31300
rect 32272 31288 32278 31340
rect 32306 31288 32312 31340
rect 32364 31328 32370 31340
rect 32401 31331 32459 31337
rect 32401 31328 32413 31331
rect 32364 31300 32413 31328
rect 32364 31288 32370 31300
rect 32401 31297 32413 31300
rect 32447 31297 32459 31331
rect 32401 31291 32459 31297
rect 33404 31331 33462 31337
rect 33404 31297 33416 31331
rect 33450 31328 33462 31331
rect 34698 31328 34704 31340
rect 33450 31300 34704 31328
rect 33450 31297 33462 31300
rect 33404 31291 33462 31297
rect 34698 31288 34704 31300
rect 34756 31288 34762 31340
rect 35710 31288 35716 31340
rect 35768 31328 35774 31340
rect 36173 31331 36231 31337
rect 36173 31328 36185 31331
rect 35768 31300 36185 31328
rect 35768 31288 35774 31300
rect 36173 31297 36185 31300
rect 36219 31297 36231 31331
rect 36173 31291 36231 31297
rect 37737 31331 37795 31337
rect 37737 31297 37749 31331
rect 37783 31328 37795 31331
rect 37826 31328 37832 31340
rect 37783 31300 37832 31328
rect 37783 31297 37795 31300
rect 37737 31291 37795 31297
rect 37826 31288 37832 31300
rect 37884 31288 37890 31340
rect 38930 31288 38936 31340
rect 38988 31328 38994 31340
rect 39025 31331 39083 31337
rect 39025 31328 39037 31331
rect 38988 31300 39037 31328
rect 38988 31288 38994 31300
rect 39025 31297 39037 31300
rect 39071 31297 39083 31331
rect 39025 31291 39083 31297
rect 39853 31331 39911 31337
rect 39853 31297 39865 31331
rect 39899 31328 39911 31331
rect 40218 31328 40224 31340
rect 39899 31300 40224 31328
rect 39899 31297 39911 31300
rect 39853 31291 39911 31297
rect 40218 31288 40224 31300
rect 40276 31288 40282 31340
rect 41877 31331 41935 31337
rect 41877 31297 41889 31331
rect 41923 31297 41935 31331
rect 42518 31328 42524 31340
rect 42479 31300 42524 31328
rect 41877 31291 41935 31297
rect 32677 31263 32735 31269
rect 32677 31229 32689 31263
rect 32723 31260 32735 31263
rect 33137 31263 33195 31269
rect 33137 31260 33149 31263
rect 32723 31232 33149 31260
rect 32723 31229 32735 31232
rect 32677 31223 32735 31229
rect 33137 31229 33149 31232
rect 33183 31229 33195 31263
rect 41892 31260 41920 31291
rect 42518 31288 42524 31300
rect 42576 31288 42582 31340
rect 42613 31331 42671 31337
rect 42613 31297 42625 31331
rect 42659 31328 42671 31331
rect 42978 31328 42984 31340
rect 42659 31300 42984 31328
rect 42659 31297 42671 31300
rect 42613 31291 42671 31297
rect 42978 31288 42984 31300
rect 43036 31328 43042 31340
rect 43036 31300 43208 31328
rect 43036 31288 43042 31300
rect 42797 31263 42855 31269
rect 42797 31260 42809 31263
rect 41892 31232 42809 31260
rect 33137 31223 33195 31229
rect 42797 31229 42809 31232
rect 42843 31229 42855 31263
rect 43180 31260 43208 31300
rect 43438 31288 43444 31340
rect 43496 31328 43502 31340
rect 43717 31331 43775 31337
rect 43717 31328 43729 31331
rect 43496 31300 43729 31328
rect 43496 31288 43502 31300
rect 43717 31297 43729 31300
rect 43763 31297 43775 31331
rect 43717 31291 43775 31297
rect 44174 31288 44180 31340
rect 44232 31328 44238 31340
rect 65812 31337 65840 31368
rect 66254 31356 66260 31368
rect 66312 31356 66318 31408
rect 44637 31331 44695 31337
rect 44637 31328 44649 31331
rect 44232 31300 44649 31328
rect 44232 31288 44238 31300
rect 44637 31297 44649 31300
rect 44683 31297 44695 31331
rect 44637 31291 44695 31297
rect 65797 31331 65855 31337
rect 65797 31297 65809 31331
rect 65843 31297 65855 31331
rect 65797 31291 65855 31297
rect 43990 31260 43996 31272
rect 43180 31232 43996 31260
rect 42797 31223 42855 31229
rect 43990 31220 43996 31232
rect 44048 31220 44054 31272
rect 65978 31260 65984 31272
rect 65939 31232 65984 31260
rect 65978 31220 65984 31232
rect 66036 31220 66042 31272
rect 67542 31260 67548 31272
rect 67503 31232 67548 31260
rect 67542 31220 67548 31232
rect 67600 31220 67606 31272
rect 35986 31192 35992 31204
rect 35544 31164 35992 31192
rect 26326 31124 26332 31136
rect 24596 31096 26332 31124
rect 26326 31084 26332 31096
rect 26384 31084 26390 31136
rect 26421 31127 26479 31133
rect 26421 31093 26433 31127
rect 26467 31124 26479 31127
rect 26510 31124 26516 31136
rect 26467 31096 26516 31124
rect 26467 31093 26479 31096
rect 26421 31087 26479 31093
rect 26510 31084 26516 31096
rect 26568 31084 26574 31136
rect 27157 31127 27215 31133
rect 27157 31093 27169 31127
rect 27203 31124 27215 31127
rect 27985 31127 28043 31133
rect 27985 31124 27997 31127
rect 27203 31096 27997 31124
rect 27203 31093 27215 31096
rect 27157 31087 27215 31093
rect 27985 31093 27997 31096
rect 28031 31124 28043 31127
rect 28074 31124 28080 31136
rect 28031 31096 28080 31124
rect 28031 31093 28043 31096
rect 27985 31087 28043 31093
rect 28074 31084 28080 31096
rect 28132 31084 28138 31136
rect 28169 31127 28227 31133
rect 28169 31093 28181 31127
rect 28215 31124 28227 31127
rect 28534 31124 28540 31136
rect 28215 31096 28540 31124
rect 28215 31093 28227 31096
rect 28169 31087 28227 31093
rect 28534 31084 28540 31096
rect 28592 31084 28598 31136
rect 31386 31124 31392 31136
rect 31347 31096 31392 31124
rect 31386 31084 31392 31096
rect 31444 31084 31450 31136
rect 33318 31084 33324 31136
rect 33376 31124 33382 31136
rect 35544 31133 35572 31164
rect 35986 31152 35992 31164
rect 36044 31152 36050 31204
rect 34517 31127 34575 31133
rect 34517 31124 34529 31127
rect 33376 31096 34529 31124
rect 33376 31084 33382 31096
rect 34517 31093 34529 31096
rect 34563 31093 34575 31127
rect 34517 31087 34575 31093
rect 35529 31127 35587 31133
rect 35529 31093 35541 31127
rect 35575 31093 35587 31127
rect 35710 31124 35716 31136
rect 35671 31096 35716 31124
rect 35529 31087 35587 31093
rect 35710 31084 35716 31096
rect 35768 31084 35774 31136
rect 36170 31124 36176 31136
rect 36131 31096 36176 31124
rect 36170 31084 36176 31096
rect 36228 31084 36234 31136
rect 37550 31124 37556 31136
rect 37511 31096 37556 31124
rect 37550 31084 37556 31096
rect 37608 31084 37614 31136
rect 39114 31084 39120 31136
rect 39172 31124 39178 31136
rect 39209 31127 39267 31133
rect 39209 31124 39221 31127
rect 39172 31096 39221 31124
rect 39172 31084 39178 31096
rect 39209 31093 39221 31096
rect 39255 31093 39267 31127
rect 43898 31124 43904 31136
rect 43859 31096 43904 31124
rect 39209 31087 39267 31093
rect 43898 31084 43904 31096
rect 43956 31084 43962 31136
rect 44450 31124 44456 31136
rect 44411 31096 44456 31124
rect 44450 31084 44456 31096
rect 44508 31084 44514 31136
rect 1104 31034 68816 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 68816 31034
rect 1104 30960 68816 30982
rect 2038 30920 2044 30932
rect 1999 30892 2044 30920
rect 2038 30880 2044 30892
rect 2096 30880 2102 30932
rect 26326 30880 26332 30932
rect 26384 30920 26390 30932
rect 26786 30920 26792 30932
rect 26384 30892 26792 30920
rect 26384 30880 26390 30892
rect 26786 30880 26792 30892
rect 26844 30920 26850 30932
rect 30466 30920 30472 30932
rect 26844 30892 30472 30920
rect 26844 30880 26850 30892
rect 30466 30880 30472 30892
rect 30524 30880 30530 30932
rect 33134 30880 33140 30932
rect 33192 30920 33198 30932
rect 33410 30920 33416 30932
rect 33192 30892 33416 30920
rect 33192 30880 33198 30892
rect 33410 30880 33416 30892
rect 33468 30880 33474 30932
rect 34698 30920 34704 30932
rect 34659 30892 34704 30920
rect 34698 30880 34704 30892
rect 34756 30880 34762 30932
rect 44174 30920 44180 30932
rect 44135 30892 44180 30920
rect 44174 30880 44180 30892
rect 44232 30880 44238 30932
rect 65978 30880 65984 30932
rect 66036 30920 66042 30932
rect 67637 30923 67695 30929
rect 67637 30920 67649 30923
rect 66036 30892 67649 30920
rect 66036 30880 66042 30892
rect 67637 30889 67649 30892
rect 67683 30889 67695 30923
rect 67637 30883 67695 30889
rect 33597 30855 33655 30861
rect 33597 30821 33609 30855
rect 33643 30821 33655 30855
rect 33597 30815 33655 30821
rect 33226 30744 33232 30796
rect 33284 30744 33290 30796
rect 1946 30716 1952 30728
rect 1859 30688 1952 30716
rect 1946 30676 1952 30688
rect 2004 30716 2010 30728
rect 3326 30716 3332 30728
rect 2004 30688 3332 30716
rect 2004 30676 2010 30688
rect 3326 30676 3332 30688
rect 3384 30676 3390 30728
rect 22462 30716 22468 30728
rect 22423 30688 22468 30716
rect 22462 30676 22468 30688
rect 22520 30676 22526 30728
rect 23198 30716 23204 30728
rect 23159 30688 23204 30716
rect 23198 30676 23204 30688
rect 23256 30676 23262 30728
rect 24578 30716 24584 30728
rect 24539 30688 24584 30716
rect 24578 30676 24584 30688
rect 24636 30676 24642 30728
rect 28534 30716 28540 30728
rect 28495 30688 28540 30716
rect 28534 30676 28540 30688
rect 28592 30676 28598 30728
rect 29549 30719 29607 30725
rect 29549 30685 29561 30719
rect 29595 30685 29607 30719
rect 31110 30716 31116 30728
rect 31071 30688 31116 30716
rect 29549 30679 29607 30685
rect 23385 30651 23443 30657
rect 23385 30617 23397 30651
rect 23431 30648 23443 30651
rect 23474 30648 23480 30660
rect 23431 30620 23480 30648
rect 23431 30617 23443 30620
rect 23385 30611 23443 30617
rect 23474 30608 23480 30620
rect 23532 30608 23538 30660
rect 29564 30648 29592 30679
rect 31110 30676 31116 30688
rect 31168 30676 31174 30728
rect 31386 30725 31392 30728
rect 31380 30716 31392 30725
rect 31347 30688 31392 30716
rect 31380 30679 31392 30688
rect 31386 30676 31392 30679
rect 31444 30676 31450 30728
rect 33244 30716 33272 30744
rect 33612 30716 33640 30815
rect 37550 30784 37556 30796
rect 37511 30756 37556 30784
rect 37550 30744 37556 30756
rect 37608 30744 37614 30796
rect 34885 30719 34943 30725
rect 34885 30716 34897 30719
rect 33244 30688 33456 30716
rect 33612 30688 34897 30716
rect 31754 30648 31760 30660
rect 29564 30620 31760 30648
rect 31754 30608 31760 30620
rect 31812 30648 31818 30660
rect 32306 30648 32312 30660
rect 31812 30620 32312 30648
rect 31812 30608 31818 30620
rect 32306 30608 32312 30620
rect 32364 30608 32370 30660
rect 33229 30651 33287 30657
rect 33229 30617 33241 30651
rect 33275 30648 33287 30651
rect 33318 30648 33324 30660
rect 33275 30620 33324 30648
rect 33275 30617 33287 30620
rect 33229 30611 33287 30617
rect 33318 30608 33324 30620
rect 33376 30608 33382 30660
rect 33428 30657 33456 30688
rect 34885 30685 34897 30688
rect 34931 30685 34943 30719
rect 34885 30679 34943 30685
rect 35529 30719 35587 30725
rect 35529 30685 35541 30719
rect 35575 30716 35587 30719
rect 36170 30716 36176 30728
rect 35575 30688 36176 30716
rect 35575 30685 35587 30688
rect 35529 30679 35587 30685
rect 36170 30676 36176 30688
rect 36228 30676 36234 30728
rect 40034 30676 40040 30728
rect 40092 30716 40098 30728
rect 40405 30719 40463 30725
rect 40405 30716 40417 30719
rect 40092 30688 40417 30716
rect 40092 30676 40098 30688
rect 40405 30685 40417 30688
rect 40451 30685 40463 30719
rect 40405 30679 40463 30685
rect 40589 30719 40647 30725
rect 40589 30685 40601 30719
rect 40635 30685 40647 30719
rect 40589 30679 40647 30685
rect 33428 30651 33487 30657
rect 33428 30620 33441 30651
rect 33429 30617 33441 30620
rect 33475 30617 33487 30651
rect 33429 30611 33487 30617
rect 35342 30608 35348 30660
rect 35400 30648 35406 30660
rect 35774 30651 35832 30657
rect 35774 30648 35786 30651
rect 35400 30620 35786 30648
rect 35400 30608 35406 30620
rect 35774 30617 35786 30620
rect 35820 30617 35832 30651
rect 35774 30611 35832 30617
rect 37820 30651 37878 30657
rect 37820 30617 37832 30651
rect 37866 30648 37878 30651
rect 38194 30648 38200 30660
rect 37866 30620 38200 30648
rect 37866 30617 37878 30620
rect 37820 30611 37878 30617
rect 38194 30608 38200 30620
rect 38252 30608 38258 30660
rect 40126 30608 40132 30660
rect 40184 30648 40190 30660
rect 40604 30648 40632 30679
rect 41138 30676 41144 30728
rect 41196 30716 41202 30728
rect 41233 30719 41291 30725
rect 41233 30716 41245 30719
rect 41196 30688 41245 30716
rect 41196 30676 41202 30688
rect 41233 30685 41245 30688
rect 41279 30685 41291 30719
rect 41233 30679 41291 30685
rect 42702 30676 42708 30728
rect 42760 30716 42766 30728
rect 42981 30719 43039 30725
rect 42981 30716 42993 30719
rect 42760 30688 42993 30716
rect 42760 30676 42766 30688
rect 42981 30685 42993 30688
rect 43027 30685 43039 30719
rect 42981 30679 43039 30685
rect 43901 30719 43959 30725
rect 43901 30685 43913 30719
rect 43947 30685 43959 30719
rect 43901 30679 43959 30685
rect 40184 30620 40632 30648
rect 43165 30651 43223 30657
rect 40184 30608 40190 30620
rect 43165 30617 43177 30651
rect 43211 30648 43223 30651
rect 43916 30648 43944 30679
rect 43990 30676 43996 30728
rect 44048 30716 44054 30728
rect 44048 30688 44093 30716
rect 44048 30676 44054 30688
rect 66806 30676 66812 30728
rect 66864 30716 66870 30728
rect 67542 30716 67548 30728
rect 66864 30688 67548 30716
rect 66864 30676 66870 30688
rect 67542 30676 67548 30688
rect 67600 30676 67606 30728
rect 45462 30648 45468 30660
rect 43211 30620 45468 30648
rect 43211 30617 43223 30620
rect 43165 30611 43223 30617
rect 45462 30608 45468 30620
rect 45520 30608 45526 30660
rect 22094 30540 22100 30592
rect 22152 30580 22158 30592
rect 22281 30583 22339 30589
rect 22281 30580 22293 30583
rect 22152 30552 22293 30580
rect 22152 30540 22158 30552
rect 22281 30549 22293 30552
rect 22327 30549 22339 30583
rect 24394 30580 24400 30592
rect 24355 30552 24400 30580
rect 22281 30543 22339 30549
rect 24394 30540 24400 30552
rect 24452 30540 24458 30592
rect 28350 30580 28356 30592
rect 28311 30552 28356 30580
rect 28350 30540 28356 30552
rect 28408 30540 28414 30592
rect 29638 30580 29644 30592
rect 29599 30552 29644 30580
rect 29638 30540 29644 30552
rect 29696 30540 29702 30592
rect 32490 30580 32496 30592
rect 32451 30552 32496 30580
rect 32490 30540 32496 30552
rect 32548 30540 32554 30592
rect 34514 30540 34520 30592
rect 34572 30580 34578 30592
rect 36909 30583 36967 30589
rect 36909 30580 36921 30583
rect 34572 30552 36921 30580
rect 34572 30540 34578 30552
rect 36909 30549 36921 30552
rect 36955 30549 36967 30583
rect 36909 30543 36967 30549
rect 38838 30540 38844 30592
rect 38896 30580 38902 30592
rect 38933 30583 38991 30589
rect 38933 30580 38945 30583
rect 38896 30552 38945 30580
rect 38896 30540 38902 30552
rect 38933 30549 38945 30552
rect 38979 30549 38991 30583
rect 40770 30580 40776 30592
rect 40731 30552 40776 30580
rect 38933 30543 38991 30549
rect 40770 30540 40776 30552
rect 40828 30540 40834 30592
rect 41414 30540 41420 30592
rect 41472 30580 41478 30592
rect 41472 30552 41517 30580
rect 41472 30540 41478 30552
rect 42978 30540 42984 30592
rect 43036 30580 43042 30592
rect 43349 30583 43407 30589
rect 43349 30580 43361 30583
rect 43036 30552 43361 30580
rect 43036 30540 43042 30552
rect 43349 30549 43361 30552
rect 43395 30549 43407 30583
rect 43349 30543 43407 30549
rect 1104 30490 68816 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 68816 30490
rect 1104 30416 68816 30438
rect 22462 30336 22468 30388
rect 22520 30376 22526 30388
rect 23017 30379 23075 30385
rect 23017 30376 23029 30379
rect 22520 30348 23029 30376
rect 22520 30336 22526 30348
rect 23017 30345 23029 30348
rect 23063 30345 23075 30379
rect 31110 30376 31116 30388
rect 31071 30348 31116 30376
rect 23017 30339 23075 30345
rect 31110 30336 31116 30348
rect 31168 30336 31174 30388
rect 32214 30336 32220 30388
rect 32272 30376 32278 30388
rect 32953 30379 33011 30385
rect 32953 30376 32965 30379
rect 32272 30348 32965 30376
rect 32272 30336 32278 30348
rect 32953 30345 32965 30348
rect 32999 30345 33011 30379
rect 34514 30376 34520 30388
rect 32953 30339 33011 30345
rect 33704 30348 34520 30376
rect 23198 30308 23204 30320
rect 22020 30280 23204 30308
rect 22020 30249 22048 30280
rect 23198 30268 23204 30280
rect 23256 30268 23262 30320
rect 23566 30308 23572 30320
rect 23308 30280 23572 30308
rect 22005 30243 22063 30249
rect 22005 30209 22017 30243
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 22833 30243 22891 30249
rect 22833 30209 22845 30243
rect 22879 30240 22891 30243
rect 23308 30240 23336 30280
rect 23566 30268 23572 30280
rect 23624 30268 23630 30320
rect 23744 30311 23802 30317
rect 23744 30277 23756 30311
rect 23790 30308 23802 30311
rect 24394 30308 24400 30320
rect 23790 30280 24400 30308
rect 23790 30277 23802 30280
rect 23744 30271 23802 30277
rect 24394 30268 24400 30280
rect 24452 30268 24458 30320
rect 28350 30268 28356 30320
rect 28408 30308 28414 30320
rect 28782 30311 28840 30317
rect 28782 30308 28794 30311
rect 28408 30280 28794 30308
rect 28408 30268 28414 30280
rect 28782 30277 28794 30280
rect 28828 30277 28840 30311
rect 28782 30271 28840 30277
rect 32122 30268 32128 30320
rect 32180 30308 32186 30320
rect 32490 30308 32496 30320
rect 32180 30280 32496 30308
rect 32180 30268 32186 30280
rect 32490 30268 32496 30280
rect 32548 30308 32554 30320
rect 32585 30311 32643 30317
rect 32585 30308 32597 30311
rect 32548 30280 32597 30308
rect 32548 30268 32554 30280
rect 32585 30277 32597 30280
rect 32631 30277 32643 30311
rect 32585 30271 32643 30277
rect 32801 30311 32859 30317
rect 32801 30277 32813 30311
rect 32847 30308 32859 30311
rect 33226 30308 33232 30320
rect 32847 30280 33232 30308
rect 32847 30277 32859 30280
rect 32801 30271 32859 30277
rect 33226 30268 33232 30280
rect 33284 30268 33290 30320
rect 23474 30240 23480 30252
rect 22879 30212 23336 30240
rect 23435 30212 23480 30240
rect 22879 30209 22891 30212
rect 22833 30203 22891 30209
rect 23474 30200 23480 30212
rect 23532 30200 23538 30252
rect 28537 30243 28595 30249
rect 28537 30209 28549 30243
rect 28583 30240 28595 30243
rect 29638 30240 29644 30252
rect 28583 30212 29644 30240
rect 28583 30209 28595 30212
rect 28537 30203 28595 30209
rect 29638 30200 29644 30212
rect 29696 30200 29702 30252
rect 31113 30243 31171 30249
rect 31113 30209 31125 30243
rect 31159 30240 31171 30243
rect 31754 30240 31760 30252
rect 31159 30212 31760 30240
rect 31159 30209 31171 30212
rect 31113 30203 31171 30209
rect 31754 30200 31760 30212
rect 31812 30200 31818 30252
rect 33318 30200 33324 30252
rect 33376 30240 33382 30252
rect 33704 30249 33732 30348
rect 34514 30336 34520 30348
rect 34572 30336 34578 30388
rect 38194 30376 38200 30388
rect 38155 30348 38200 30376
rect 38194 30336 38200 30348
rect 38252 30336 38258 30388
rect 40034 30336 40040 30388
rect 40092 30376 40098 30388
rect 41877 30379 41935 30385
rect 41877 30376 41889 30379
rect 40092 30348 41889 30376
rect 40092 30336 40098 30348
rect 41877 30345 41889 30348
rect 41923 30345 41935 30379
rect 45462 30376 45468 30388
rect 45423 30348 45468 30376
rect 41877 30339 41935 30345
rect 45462 30336 45468 30348
rect 45520 30336 45526 30388
rect 36541 30311 36599 30317
rect 36541 30277 36553 30311
rect 36587 30308 36599 30311
rect 37366 30308 37372 30320
rect 36587 30280 37372 30308
rect 36587 30277 36599 30280
rect 36541 30271 36599 30277
rect 37366 30268 37372 30280
rect 37424 30308 37430 30320
rect 37461 30311 37519 30317
rect 37461 30308 37473 30311
rect 37424 30280 37473 30308
rect 37424 30268 37430 30280
rect 37461 30277 37473 30280
rect 37507 30277 37519 30311
rect 41414 30308 41420 30320
rect 37461 30271 37519 30277
rect 40512 30280 41420 30308
rect 33505 30243 33563 30249
rect 33505 30240 33517 30243
rect 33376 30212 33517 30240
rect 33376 30200 33382 30212
rect 33505 30209 33517 30212
rect 33551 30209 33563 30243
rect 33505 30203 33563 30209
rect 33689 30243 33747 30249
rect 33689 30209 33701 30243
rect 33735 30209 33747 30243
rect 33689 30203 33747 30209
rect 35345 30243 35403 30249
rect 35345 30209 35357 30243
rect 35391 30240 35403 30243
rect 36357 30243 36415 30249
rect 36357 30240 36369 30243
rect 35391 30212 36369 30240
rect 35391 30209 35403 30212
rect 35345 30203 35403 30209
rect 36357 30209 36369 30212
rect 36403 30209 36415 30243
rect 36357 30203 36415 30209
rect 37277 30243 37335 30249
rect 37277 30209 37289 30243
rect 37323 30209 37335 30243
rect 38378 30240 38384 30252
rect 38339 30212 38384 30240
rect 37277 30203 37335 30209
rect 1854 30172 1860 30184
rect 1815 30144 1860 30172
rect 1854 30132 1860 30144
rect 1912 30132 1918 30184
rect 2041 30175 2099 30181
rect 2041 30141 2053 30175
rect 2087 30172 2099 30175
rect 2774 30172 2780 30184
rect 2087 30144 2780 30172
rect 2087 30141 2099 30144
rect 2041 30135 2099 30141
rect 2774 30132 2780 30144
rect 2832 30132 2838 30184
rect 2866 30132 2872 30184
rect 2924 30172 2930 30184
rect 22649 30175 22707 30181
rect 2924 30144 2969 30172
rect 2924 30132 2930 30144
rect 22649 30141 22661 30175
rect 22695 30172 22707 30175
rect 23198 30172 23204 30184
rect 22695 30144 23204 30172
rect 22695 30141 22707 30144
rect 22649 30135 22707 30141
rect 23198 30132 23204 30144
rect 23256 30132 23262 30184
rect 34054 30132 34060 30184
rect 34112 30172 34118 30184
rect 34425 30175 34483 30181
rect 34425 30172 34437 30175
rect 34112 30144 34437 30172
rect 34112 30132 34118 30144
rect 34425 30141 34437 30144
rect 34471 30141 34483 30175
rect 34425 30135 34483 30141
rect 34514 30132 34520 30184
rect 34572 30181 34578 30184
rect 34572 30175 34600 30181
rect 34588 30141 34600 30175
rect 34572 30135 34600 30141
rect 34572 30132 34578 30135
rect 34698 30132 34704 30184
rect 34756 30172 34762 30184
rect 34882 30172 34888 30184
rect 34756 30144 34888 30172
rect 34756 30132 34762 30144
rect 34882 30132 34888 30144
rect 34940 30132 34946 30184
rect 37292 30172 37320 30203
rect 38378 30200 38384 30212
rect 38436 30200 38442 30252
rect 39114 30240 39120 30252
rect 39075 30212 39120 30240
rect 39114 30200 39120 30212
rect 39172 30200 39178 30252
rect 39301 30243 39359 30249
rect 39301 30209 39313 30243
rect 39347 30240 39359 30243
rect 39482 30240 39488 30252
rect 39347 30212 39488 30240
rect 39347 30209 39359 30212
rect 39301 30203 39359 30209
rect 39482 30200 39488 30212
rect 39540 30200 39546 30252
rect 40512 30249 40540 30280
rect 41414 30268 41420 30280
rect 41472 30268 41478 30320
rect 43254 30308 43260 30320
rect 43180 30280 43260 30308
rect 40497 30243 40555 30249
rect 40497 30209 40509 30243
rect 40543 30209 40555 30243
rect 40497 30203 40555 30209
rect 40586 30200 40592 30252
rect 40644 30240 40650 30252
rect 40753 30243 40811 30249
rect 40753 30240 40765 30243
rect 40644 30212 40765 30240
rect 40644 30200 40650 30212
rect 40753 30209 40765 30212
rect 40799 30209 40811 30243
rect 42978 30240 42984 30252
rect 42939 30212 42984 30240
rect 40753 30203 40811 30209
rect 42978 30200 42984 30212
rect 43036 30200 43042 30252
rect 43180 30249 43208 30280
rect 43254 30268 43260 30280
rect 43312 30268 43318 30320
rect 44352 30311 44410 30317
rect 44352 30277 44364 30311
rect 44398 30308 44410 30311
rect 44450 30308 44456 30320
rect 44398 30280 44456 30308
rect 44398 30277 44410 30280
rect 44352 30271 44410 30277
rect 44450 30268 44456 30280
rect 44508 30268 44514 30320
rect 49602 30268 49608 30320
rect 49660 30308 49666 30320
rect 66162 30308 66168 30320
rect 49660 30280 66168 30308
rect 49660 30268 49666 30280
rect 66162 30268 66168 30280
rect 66220 30268 66226 30320
rect 43165 30243 43223 30249
rect 43165 30209 43177 30243
rect 43211 30209 43223 30243
rect 43165 30203 43223 30209
rect 43898 30200 43904 30252
rect 43956 30240 43962 30252
rect 44085 30243 44143 30249
rect 44085 30240 44097 30243
rect 43956 30212 44097 30240
rect 43956 30200 43962 30212
rect 44085 30209 44097 30212
rect 44131 30209 44143 30243
rect 44085 30203 44143 30209
rect 35084 30144 37320 30172
rect 37645 30175 37703 30181
rect 24486 30064 24492 30116
rect 24544 30104 24550 30116
rect 28074 30104 28080 30116
rect 24544 30076 28080 30104
rect 24544 30064 24550 30076
rect 28074 30064 28080 30076
rect 28132 30064 28138 30116
rect 29822 30064 29828 30116
rect 29880 30104 29886 30116
rect 32674 30104 32680 30116
rect 29880 30076 32680 30104
rect 29880 30064 29886 30076
rect 32674 30064 32680 30076
rect 32732 30064 32738 30116
rect 33410 30104 33416 30116
rect 32784 30076 33416 30104
rect 21818 29996 21824 30048
rect 21876 30036 21882 30048
rect 21913 30039 21971 30045
rect 21913 30036 21925 30039
rect 21876 30008 21925 30036
rect 21876 29996 21882 30008
rect 21913 30005 21925 30008
rect 21959 30005 21971 30039
rect 21913 29999 21971 30005
rect 24394 29996 24400 30048
rect 24452 30036 24458 30048
rect 24857 30039 24915 30045
rect 24857 30036 24869 30039
rect 24452 30008 24869 30036
rect 24452 29996 24458 30008
rect 24857 30005 24869 30008
rect 24903 30036 24915 30039
rect 27338 30036 27344 30048
rect 24903 30008 27344 30036
rect 24903 30005 24915 30008
rect 24857 29999 24915 30005
rect 27338 29996 27344 30008
rect 27396 29996 27402 30048
rect 27798 29996 27804 30048
rect 27856 30036 27862 30048
rect 32784 30045 32812 30076
rect 33410 30064 33416 30076
rect 33468 30064 33474 30116
rect 34146 30104 34152 30116
rect 34107 30076 34152 30104
rect 34146 30064 34152 30076
rect 34204 30064 34210 30116
rect 29917 30039 29975 30045
rect 29917 30036 29929 30039
rect 27856 30008 29929 30036
rect 27856 29996 27862 30008
rect 29917 30005 29929 30008
rect 29963 30005 29975 30039
rect 29917 29999 29975 30005
rect 32769 30039 32827 30045
rect 32769 30005 32781 30039
rect 32815 30005 32827 30039
rect 32769 29999 32827 30005
rect 34422 29996 34428 30048
rect 34480 30036 34486 30048
rect 35084 30036 35112 30144
rect 37645 30141 37657 30175
rect 37691 30172 37703 30175
rect 39209 30175 39267 30181
rect 39209 30172 39221 30175
rect 37691 30144 39221 30172
rect 37691 30141 37703 30144
rect 37645 30135 37703 30141
rect 39209 30141 39221 30144
rect 39255 30141 39267 30175
rect 39209 30135 39267 30141
rect 39393 30175 39451 30181
rect 39393 30141 39405 30175
rect 39439 30172 39451 30175
rect 40310 30172 40316 30184
rect 39439 30144 40316 30172
rect 39439 30141 39451 30144
rect 39393 30135 39451 30141
rect 40310 30132 40316 30144
rect 40368 30132 40374 30184
rect 43073 30175 43131 30181
rect 43073 30141 43085 30175
rect 43119 30141 43131 30175
rect 43073 30135 43131 30141
rect 43257 30175 43315 30181
rect 43257 30141 43269 30175
rect 43303 30172 43315 30175
rect 43622 30172 43628 30184
rect 43303 30144 43628 30172
rect 43303 30141 43315 30144
rect 43257 30135 43315 30141
rect 36725 30107 36783 30113
rect 36725 30073 36737 30107
rect 36771 30104 36783 30107
rect 43088 30104 43116 30135
rect 43622 30132 43628 30144
rect 43680 30132 43686 30184
rect 36771 30076 39068 30104
rect 36771 30073 36783 30076
rect 36725 30067 36783 30073
rect 38930 30036 38936 30048
rect 34480 30008 35112 30036
rect 38891 30008 38936 30036
rect 34480 29996 34486 30008
rect 38930 29996 38936 30008
rect 38988 29996 38994 30048
rect 39040 30036 39068 30076
rect 42260 30076 43116 30104
rect 42260 30036 42288 30076
rect 39040 30008 42288 30036
rect 42797 30039 42855 30045
rect 42797 30005 42809 30039
rect 42843 30036 42855 30039
rect 43254 30036 43260 30048
rect 42843 30008 43260 30036
rect 42843 30005 42855 30008
rect 42797 29999 42855 30005
rect 43254 29996 43260 30008
rect 43312 29996 43318 30048
rect 1104 29946 68816 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 68816 29946
rect 1104 29872 68816 29894
rect 1854 29792 1860 29844
rect 1912 29832 1918 29844
rect 2041 29835 2099 29841
rect 2041 29832 2053 29835
rect 1912 29804 2053 29832
rect 1912 29792 1918 29804
rect 2041 29801 2053 29804
rect 2087 29801 2099 29835
rect 2774 29832 2780 29844
rect 2735 29804 2780 29832
rect 2041 29795 2099 29801
rect 2774 29792 2780 29804
rect 2832 29792 2838 29844
rect 23198 29832 23204 29844
rect 23111 29804 23204 29832
rect 23198 29792 23204 29804
rect 23256 29832 23262 29844
rect 24486 29832 24492 29844
rect 23256 29804 24492 29832
rect 23256 29792 23262 29804
rect 24486 29792 24492 29804
rect 24544 29792 24550 29844
rect 24578 29792 24584 29844
rect 24636 29832 24642 29844
rect 24765 29835 24823 29841
rect 24765 29832 24777 29835
rect 24636 29804 24777 29832
rect 24636 29792 24642 29804
rect 24765 29801 24777 29804
rect 24811 29801 24823 29835
rect 27706 29832 27712 29844
rect 24765 29795 24823 29801
rect 27080 29804 27712 29832
rect 27080 29773 27108 29804
rect 27706 29792 27712 29804
rect 27764 29792 27770 29844
rect 28261 29835 28319 29841
rect 28261 29801 28273 29835
rect 28307 29832 28319 29835
rect 34422 29832 34428 29844
rect 28307 29804 34428 29832
rect 28307 29801 28319 29804
rect 28261 29795 28319 29801
rect 34422 29792 34428 29804
rect 34480 29792 34486 29844
rect 35342 29832 35348 29844
rect 35303 29804 35348 29832
rect 35342 29792 35348 29804
rect 35400 29792 35406 29844
rect 38378 29792 38384 29844
rect 38436 29832 38442 29844
rect 39117 29835 39175 29841
rect 39117 29832 39129 29835
rect 38436 29804 39129 29832
rect 38436 29792 38442 29804
rect 39117 29801 39129 29804
rect 39163 29801 39175 29835
rect 39117 29795 39175 29801
rect 27065 29767 27123 29773
rect 26206 29736 26648 29764
rect 21818 29696 21824 29708
rect 21779 29668 21824 29696
rect 21818 29656 21824 29668
rect 21876 29656 21882 29708
rect 24394 29696 24400 29708
rect 24355 29668 24400 29696
rect 24394 29656 24400 29668
rect 24452 29656 24458 29708
rect 2685 29631 2743 29637
rect 2685 29597 2697 29631
rect 2731 29628 2743 29631
rect 4798 29628 4804 29640
rect 2731 29600 4804 29628
rect 2731 29597 2743 29600
rect 2685 29591 2743 29597
rect 4798 29588 4804 29600
rect 4856 29588 4862 29640
rect 22094 29637 22100 29640
rect 22088 29628 22100 29637
rect 22055 29600 22100 29628
rect 22088 29591 22100 29600
rect 22094 29588 22100 29591
rect 22152 29588 22158 29640
rect 23566 29588 23572 29640
rect 23624 29628 23630 29640
rect 24581 29631 24639 29637
rect 24581 29628 24593 29631
rect 23624 29600 24593 29628
rect 23624 29588 23630 29600
rect 24581 29597 24593 29600
rect 24627 29597 24639 29631
rect 24581 29591 24639 29597
rect 25409 29631 25467 29637
rect 25409 29597 25421 29631
rect 25455 29628 25467 29631
rect 25682 29628 25688 29640
rect 25455 29600 25688 29628
rect 25455 29597 25467 29600
rect 25409 29591 25467 29597
rect 25682 29588 25688 29600
rect 25740 29588 25746 29640
rect 25222 29492 25228 29504
rect 25183 29464 25228 29492
rect 25222 29452 25228 29464
rect 25280 29452 25286 29504
rect 26050 29452 26056 29504
rect 26108 29492 26114 29504
rect 26206 29492 26234 29736
rect 26421 29699 26479 29705
rect 26421 29665 26433 29699
rect 26467 29696 26479 29699
rect 26510 29696 26516 29708
rect 26467 29668 26516 29696
rect 26467 29665 26479 29668
rect 26421 29659 26479 29665
rect 26510 29656 26516 29668
rect 26568 29656 26574 29708
rect 26620 29696 26648 29736
rect 27065 29733 27077 29767
rect 27111 29733 27123 29767
rect 27065 29727 27123 29733
rect 31113 29767 31171 29773
rect 31113 29733 31125 29767
rect 31159 29733 31171 29767
rect 31113 29727 31171 29733
rect 27458 29699 27516 29705
rect 27458 29696 27470 29699
rect 26620 29668 27470 29696
rect 27458 29665 27470 29668
rect 27504 29665 27516 29699
rect 27458 29659 27516 29665
rect 27617 29699 27675 29705
rect 27617 29665 27629 29699
rect 27663 29696 27675 29699
rect 31128 29696 31156 29727
rect 32674 29724 32680 29776
rect 32732 29764 32738 29776
rect 34698 29764 34704 29776
rect 32732 29736 34704 29764
rect 32732 29724 32738 29736
rect 34698 29724 34704 29736
rect 34756 29724 34762 29776
rect 31573 29699 31631 29705
rect 31573 29696 31585 29699
rect 27663 29668 29868 29696
rect 31128 29668 31585 29696
rect 27663 29665 27675 29668
rect 27617 29659 27675 29665
rect 29840 29640 29868 29668
rect 31573 29665 31585 29668
rect 31619 29696 31631 29699
rect 34514 29696 34520 29708
rect 31619 29668 34520 29696
rect 31619 29665 31631 29668
rect 31573 29659 31631 29665
rect 34514 29656 34520 29668
rect 34572 29656 34578 29708
rect 37185 29699 37243 29705
rect 37185 29665 37197 29699
rect 37231 29696 37243 29699
rect 40957 29699 41015 29705
rect 40957 29696 40969 29699
rect 37231 29668 40969 29696
rect 37231 29665 37243 29668
rect 37185 29659 37243 29665
rect 40957 29665 40969 29668
rect 41003 29665 41015 29699
rect 40957 29659 41015 29665
rect 41049 29699 41107 29705
rect 41049 29665 41061 29699
rect 41095 29696 41107 29699
rect 43162 29696 43168 29708
rect 41095 29668 43168 29696
rect 41095 29665 41107 29668
rect 41049 29659 41107 29665
rect 43162 29656 43168 29668
rect 43220 29656 43226 29708
rect 26605 29631 26663 29637
rect 26605 29597 26617 29631
rect 26651 29597 26663 29631
rect 26605 29591 26663 29597
rect 26108 29464 26234 29492
rect 26620 29492 26648 29591
rect 27338 29588 27344 29640
rect 27396 29628 27402 29640
rect 27396 29600 27441 29628
rect 27396 29588 27402 29600
rect 29638 29588 29644 29640
rect 29696 29628 29702 29640
rect 29733 29631 29791 29637
rect 29733 29628 29745 29631
rect 29696 29600 29745 29628
rect 29696 29588 29702 29600
rect 29733 29597 29745 29600
rect 29779 29597 29791 29631
rect 29733 29591 29791 29597
rect 29822 29588 29828 29640
rect 29880 29588 29886 29640
rect 31757 29631 31815 29637
rect 31757 29597 31769 29631
rect 31803 29628 31815 29631
rect 31846 29628 31852 29640
rect 31803 29600 31852 29628
rect 31803 29597 31815 29600
rect 31757 29591 31815 29597
rect 31846 29588 31852 29600
rect 31904 29588 31910 29640
rect 35529 29631 35587 29637
rect 35529 29597 35541 29631
rect 35575 29628 35587 29631
rect 35710 29628 35716 29640
rect 35575 29600 35716 29628
rect 35575 29597 35587 29600
rect 35529 29591 35587 29597
rect 35710 29588 35716 29600
rect 35768 29588 35774 29640
rect 37001 29631 37059 29637
rect 37001 29597 37013 29631
rect 37047 29628 37059 29631
rect 37366 29628 37372 29640
rect 37047 29600 37372 29628
rect 37047 29597 37059 29600
rect 37001 29591 37059 29597
rect 37366 29588 37372 29600
rect 37424 29588 37430 29640
rect 38838 29628 38844 29640
rect 38799 29600 38844 29628
rect 38838 29588 38844 29600
rect 38896 29588 38902 29640
rect 38933 29631 38991 29637
rect 38933 29597 38945 29631
rect 38979 29597 38991 29631
rect 38933 29591 38991 29597
rect 30000 29563 30058 29569
rect 30000 29529 30012 29563
rect 30046 29560 30058 29563
rect 30282 29560 30288 29572
rect 30046 29532 30288 29560
rect 30046 29529 30058 29532
rect 30000 29523 30058 29529
rect 30282 29520 30288 29532
rect 30340 29520 30346 29572
rect 36817 29563 36875 29569
rect 36817 29560 36829 29563
rect 31036 29532 36829 29560
rect 27614 29492 27620 29504
rect 26620 29464 27620 29492
rect 26108 29452 26114 29464
rect 27614 29452 27620 29464
rect 27672 29452 27678 29504
rect 28994 29452 29000 29504
rect 29052 29492 29058 29504
rect 31036 29492 31064 29532
rect 36817 29529 36829 29532
rect 36863 29529 36875 29563
rect 38948 29560 38976 29591
rect 39206 29588 39212 29640
rect 39264 29628 39270 29640
rect 39853 29631 39911 29637
rect 39853 29628 39865 29631
rect 39264 29600 39865 29628
rect 39264 29588 39270 29600
rect 39853 29597 39865 29600
rect 39899 29597 39911 29631
rect 40034 29628 40040 29640
rect 39995 29600 40040 29628
rect 39853 29591 39911 29597
rect 40034 29588 40040 29600
rect 40092 29588 40098 29640
rect 40221 29631 40279 29637
rect 40221 29597 40233 29631
rect 40267 29628 40279 29631
rect 40865 29631 40923 29637
rect 40865 29628 40877 29631
rect 40267 29600 40877 29628
rect 40267 29597 40279 29600
rect 40221 29591 40279 29597
rect 40865 29597 40877 29600
rect 40911 29597 40923 29631
rect 40865 29591 40923 29597
rect 41141 29631 41199 29637
rect 41141 29597 41153 29631
rect 41187 29628 41199 29631
rect 43622 29628 43628 29640
rect 41187 29600 43628 29628
rect 41187 29597 41199 29600
rect 41141 29591 41199 29597
rect 40126 29560 40132 29572
rect 38948 29532 40132 29560
rect 36817 29523 36875 29529
rect 40126 29520 40132 29532
rect 40184 29520 40190 29572
rect 40310 29520 40316 29572
rect 40368 29560 40374 29572
rect 41156 29560 41184 29591
rect 43622 29588 43628 29600
rect 43680 29588 43686 29640
rect 45005 29631 45063 29637
rect 45005 29597 45017 29631
rect 45051 29628 45063 29631
rect 46842 29628 46848 29640
rect 45051 29600 46848 29628
rect 45051 29597 45063 29600
rect 45005 29591 45063 29597
rect 46842 29588 46848 29600
rect 46900 29588 46906 29640
rect 40368 29532 41184 29560
rect 40368 29520 40374 29532
rect 31938 29492 31944 29504
rect 29052 29464 31064 29492
rect 31899 29464 31944 29492
rect 29052 29452 29058 29464
rect 31938 29452 31944 29464
rect 31996 29452 32002 29504
rect 38930 29452 38936 29504
rect 38988 29492 38994 29504
rect 39482 29492 39488 29504
rect 38988 29464 39488 29492
rect 38988 29452 38994 29464
rect 39482 29452 39488 29464
rect 39540 29452 39546 29504
rect 40678 29492 40684 29504
rect 40639 29464 40684 29492
rect 40678 29452 40684 29464
rect 40736 29452 40742 29504
rect 44266 29452 44272 29504
rect 44324 29492 44330 29504
rect 45097 29495 45155 29501
rect 45097 29492 45109 29495
rect 44324 29464 45109 29492
rect 44324 29452 44330 29464
rect 45097 29461 45109 29464
rect 45143 29461 45155 29495
rect 45097 29455 45155 29461
rect 1104 29402 68816 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 68816 29402
rect 1104 29328 68816 29350
rect 27798 29288 27804 29300
rect 27172 29260 27804 29288
rect 24940 29223 24998 29229
rect 24940 29189 24952 29223
rect 24986 29220 24998 29223
rect 25222 29220 25228 29232
rect 24986 29192 25228 29220
rect 24986 29189 24998 29192
rect 24940 29183 24998 29189
rect 25222 29180 25228 29192
rect 25280 29180 25286 29232
rect 27172 29161 27200 29260
rect 27798 29248 27804 29260
rect 27856 29248 27862 29300
rect 27890 29248 27896 29300
rect 27948 29288 27954 29300
rect 28994 29288 29000 29300
rect 27948 29260 28856 29288
rect 28955 29260 29000 29288
rect 27948 29248 27954 29260
rect 28828 29220 28856 29260
rect 28994 29248 29000 29260
rect 29052 29248 29058 29300
rect 29638 29288 29644 29300
rect 29599 29260 29644 29288
rect 29638 29248 29644 29260
rect 29696 29248 29702 29300
rect 30282 29288 30288 29300
rect 30243 29260 30288 29288
rect 30282 29248 30288 29260
rect 30340 29248 30346 29300
rect 33962 29288 33968 29300
rect 32324 29260 33824 29288
rect 33923 29260 33968 29288
rect 28828 29192 30420 29220
rect 27157 29155 27215 29161
rect 27157 29121 27169 29155
rect 27203 29121 27215 29155
rect 27157 29115 27215 29121
rect 28074 29112 28080 29164
rect 28132 29152 28138 29164
rect 29638 29152 29644 29164
rect 28132 29124 28177 29152
rect 29599 29124 29644 29152
rect 28132 29112 28138 29124
rect 29638 29112 29644 29124
rect 29696 29112 29702 29164
rect 24670 29084 24676 29096
rect 24631 29056 24676 29084
rect 24670 29044 24676 29056
rect 24728 29044 24734 29096
rect 27341 29087 27399 29093
rect 27341 29053 27353 29087
rect 27387 29053 27399 29087
rect 27341 29047 27399 29053
rect 27356 29016 27384 29047
rect 27430 29044 27436 29096
rect 27488 29084 27494 29096
rect 28194 29087 28252 29093
rect 28194 29084 28206 29087
rect 27488 29056 28206 29084
rect 27488 29044 27494 29056
rect 28194 29053 28206 29056
rect 28240 29053 28252 29087
rect 28194 29047 28252 29053
rect 28353 29087 28411 29093
rect 28353 29053 28365 29087
rect 28399 29084 28411 29087
rect 29822 29084 29828 29096
rect 28399 29056 29828 29084
rect 28399 29053 28411 29056
rect 28353 29047 28411 29053
rect 29822 29044 29828 29056
rect 29880 29044 29886 29096
rect 27356 28988 27752 29016
rect 26050 28948 26056 28960
rect 26011 28920 26056 28948
rect 26050 28908 26056 28920
rect 26108 28908 26114 28960
rect 27724 28948 27752 28988
rect 27798 28976 27804 29028
rect 27856 29016 27862 29028
rect 30392 29016 30420 29192
rect 30469 29155 30527 29161
rect 30469 29121 30481 29155
rect 30515 29152 30527 29155
rect 31938 29152 31944 29164
rect 30515 29124 31944 29152
rect 30515 29121 30527 29124
rect 30469 29115 30527 29121
rect 31938 29112 31944 29124
rect 31996 29112 32002 29164
rect 32122 29152 32128 29164
rect 32083 29124 32128 29152
rect 32122 29112 32128 29124
rect 32180 29112 32186 29164
rect 32324 29161 32352 29260
rect 33796 29220 33824 29260
rect 33962 29248 33968 29260
rect 34020 29248 34026 29300
rect 35250 29248 35256 29300
rect 35308 29297 35314 29300
rect 35308 29291 35327 29297
rect 35315 29257 35327 29291
rect 35308 29251 35327 29257
rect 35437 29291 35495 29297
rect 35437 29257 35449 29291
rect 35483 29257 35495 29291
rect 40586 29288 40592 29300
rect 40547 29260 40592 29288
rect 35437 29251 35495 29257
rect 35308 29248 35314 29251
rect 35069 29223 35127 29229
rect 35069 29220 35081 29223
rect 33796 29192 35081 29220
rect 35069 29189 35081 29192
rect 35115 29189 35127 29223
rect 35069 29183 35127 29189
rect 32309 29155 32367 29161
rect 32309 29121 32321 29155
rect 32355 29121 32367 29155
rect 32309 29115 32367 29121
rect 32490 29044 32496 29096
rect 32548 29084 32554 29096
rect 33045 29087 33103 29093
rect 33045 29084 33057 29087
rect 32548 29056 33057 29084
rect 32548 29044 32554 29056
rect 33045 29053 33057 29056
rect 33091 29053 33103 29087
rect 33045 29047 33103 29053
rect 33134 29044 33140 29096
rect 33192 29093 33198 29096
rect 33192 29087 33220 29093
rect 33208 29053 33220 29087
rect 33192 29047 33220 29053
rect 33321 29087 33379 29093
rect 33321 29053 33333 29087
rect 33367 29084 33379 29087
rect 34698 29084 34704 29096
rect 33367 29056 34704 29084
rect 33367 29053 33379 29056
rect 33321 29047 33379 29053
rect 33192 29044 33198 29047
rect 34698 29044 34704 29056
rect 34756 29044 34762 29096
rect 35084 29084 35112 29183
rect 35452 29152 35480 29251
rect 40586 29248 40592 29260
rect 40644 29248 40650 29300
rect 44358 29288 44364 29300
rect 43180 29260 44364 29288
rect 38102 29180 38108 29232
rect 38160 29220 38166 29232
rect 38160 29192 38424 29220
rect 38160 29180 38166 29192
rect 36081 29155 36139 29161
rect 36081 29152 36093 29155
rect 35452 29124 36093 29152
rect 36081 29121 36093 29124
rect 36127 29121 36139 29155
rect 38194 29152 38200 29164
rect 38155 29124 38200 29152
rect 36081 29115 36139 29121
rect 38194 29112 38200 29124
rect 38252 29112 38258 29164
rect 38396 29161 38424 29192
rect 38580 29192 41414 29220
rect 38580 29161 38608 29192
rect 38289 29155 38347 29161
rect 38289 29121 38301 29155
rect 38335 29121 38347 29155
rect 38289 29115 38347 29121
rect 38381 29155 38439 29161
rect 38381 29121 38393 29155
rect 38427 29121 38439 29155
rect 38381 29115 38439 29121
rect 38565 29155 38623 29161
rect 38565 29121 38577 29155
rect 38611 29121 38623 29155
rect 39298 29152 39304 29164
rect 39259 29124 39304 29152
rect 38565 29115 38623 29121
rect 36538 29084 36544 29096
rect 35084 29056 36544 29084
rect 36538 29044 36544 29056
rect 36596 29044 36602 29096
rect 38304 29084 38332 29115
rect 39298 29112 39304 29124
rect 39356 29112 39362 29164
rect 39393 29155 39451 29161
rect 39393 29121 39405 29155
rect 39439 29121 39451 29155
rect 39393 29115 39451 29121
rect 39408 29084 39436 29115
rect 39482 29112 39488 29164
rect 39540 29152 39546 29164
rect 39684 29161 39712 29192
rect 39669 29155 39727 29161
rect 39540 29124 39585 29152
rect 39540 29112 39546 29124
rect 39669 29121 39681 29155
rect 39715 29121 39727 29155
rect 39669 29115 39727 29121
rect 40218 29112 40224 29164
rect 40276 29112 40282 29164
rect 40770 29152 40776 29164
rect 40731 29124 40776 29152
rect 40770 29112 40776 29124
rect 40828 29112 40834 29164
rect 40236 29084 40264 29112
rect 38304 29056 40264 29084
rect 32769 29019 32827 29025
rect 32769 29016 32781 29019
rect 27856 28988 27901 29016
rect 30392 28988 32781 29016
rect 27856 28976 27862 28988
rect 32769 28985 32781 28988
rect 32815 29016 32827 29019
rect 34146 29016 34152 29028
rect 32815 28988 32904 29016
rect 32815 28985 32827 28988
rect 32769 28979 32827 28985
rect 28810 28948 28816 28960
rect 27724 28920 28816 28948
rect 28810 28908 28816 28920
rect 28868 28908 28874 28960
rect 32876 28948 32904 28988
rect 33704 28988 34152 29016
rect 33704 28948 33732 28988
rect 34146 28976 34152 28988
rect 34204 28976 34210 29028
rect 35986 29016 35992 29028
rect 35728 28988 35992 29016
rect 32876 28920 33732 28948
rect 34698 28908 34704 28960
rect 34756 28948 34762 28960
rect 35253 28951 35311 28957
rect 35253 28948 35265 28951
rect 34756 28920 35265 28948
rect 34756 28908 34762 28920
rect 35253 28917 35265 28920
rect 35299 28948 35311 28951
rect 35728 28948 35756 28988
rect 35986 28976 35992 28988
rect 36044 28976 36050 29028
rect 39298 28976 39304 29028
rect 39356 29016 39362 29028
rect 40218 29016 40224 29028
rect 39356 28988 40224 29016
rect 39356 28976 39362 28988
rect 40218 28976 40224 28988
rect 40276 28976 40282 29028
rect 41386 29016 41414 29192
rect 43180 29161 43208 29260
rect 44358 29248 44364 29260
rect 44416 29248 44422 29300
rect 44266 29220 44272 29232
rect 44227 29192 44272 29220
rect 44266 29180 44272 29192
rect 44324 29180 44330 29232
rect 43073 29155 43131 29161
rect 43073 29121 43085 29155
rect 43119 29121 43131 29155
rect 43073 29115 43131 29121
rect 43165 29155 43223 29161
rect 43165 29121 43177 29155
rect 43211 29121 43223 29155
rect 43165 29115 43223 29121
rect 43088 29084 43116 29115
rect 43254 29112 43260 29164
rect 43312 29152 43318 29164
rect 43441 29155 43499 29161
rect 43312 29124 43357 29152
rect 43312 29112 43318 29124
rect 43441 29121 43453 29155
rect 43487 29152 43499 29155
rect 43714 29152 43720 29164
rect 43487 29124 43720 29152
rect 43487 29121 43499 29124
rect 43441 29115 43499 29121
rect 43714 29112 43720 29124
rect 43772 29112 43778 29164
rect 44085 29087 44143 29093
rect 44085 29084 44097 29087
rect 43088 29056 44097 29084
rect 44085 29053 44097 29056
rect 44131 29053 44143 29087
rect 45922 29084 45928 29096
rect 45883 29056 45928 29084
rect 44085 29047 44143 29053
rect 41506 29016 41512 29028
rect 41386 28988 41512 29016
rect 41506 28976 41512 28988
rect 41564 29016 41570 29028
rect 43714 29016 43720 29028
rect 41564 28988 43720 29016
rect 41564 28976 41570 28988
rect 43714 28976 43720 28988
rect 43772 28976 43778 29028
rect 44100 29016 44128 29047
rect 45922 29044 45928 29056
rect 45980 29044 45986 29096
rect 44174 29016 44180 29028
rect 44100 28988 44180 29016
rect 44174 28976 44180 28988
rect 44232 28976 44238 29028
rect 35894 28948 35900 28960
rect 35299 28920 35756 28948
rect 35855 28920 35900 28948
rect 35299 28917 35311 28920
rect 35253 28911 35311 28917
rect 35894 28908 35900 28920
rect 35952 28908 35958 28960
rect 37918 28948 37924 28960
rect 37879 28920 37924 28948
rect 37918 28908 37924 28920
rect 37976 28908 37982 28960
rect 39025 28951 39083 28957
rect 39025 28917 39037 28951
rect 39071 28948 39083 28951
rect 39114 28948 39120 28960
rect 39071 28920 39120 28948
rect 39071 28917 39083 28920
rect 39025 28911 39083 28917
rect 39114 28908 39120 28920
rect 39172 28908 39178 28960
rect 42797 28951 42855 28957
rect 42797 28917 42809 28951
rect 42843 28948 42855 28951
rect 42886 28948 42892 28960
rect 42843 28920 42892 28948
rect 42843 28917 42855 28920
rect 42797 28911 42855 28917
rect 42886 28908 42892 28920
rect 42944 28908 42950 28960
rect 1104 28858 68816 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 68816 28858
rect 1104 28784 68816 28806
rect 24670 28704 24676 28756
rect 24728 28744 24734 28756
rect 24765 28747 24823 28753
rect 24765 28744 24777 28747
rect 24728 28716 24777 28744
rect 24728 28704 24734 28716
rect 24765 28713 24777 28716
rect 24811 28713 24823 28747
rect 25682 28744 25688 28756
rect 25643 28716 25688 28744
rect 24765 28707 24823 28713
rect 25682 28704 25688 28716
rect 25740 28704 25746 28756
rect 29086 28704 29092 28756
rect 29144 28744 29150 28756
rect 34698 28744 34704 28756
rect 29144 28716 34704 28744
rect 29144 28704 29150 28716
rect 34698 28704 34704 28716
rect 34756 28704 34762 28756
rect 36538 28744 36544 28756
rect 36499 28716 36544 28744
rect 36538 28704 36544 28716
rect 36596 28704 36602 28756
rect 44174 28744 44180 28756
rect 44135 28716 44180 28744
rect 44174 28704 44180 28716
rect 44232 28704 44238 28756
rect 25317 28611 25375 28617
rect 25317 28577 25329 28611
rect 25363 28608 25375 28611
rect 26050 28608 26056 28620
rect 25363 28580 26056 28608
rect 25363 28577 25375 28580
rect 25317 28571 25375 28577
rect 26050 28568 26056 28580
rect 26108 28568 26114 28620
rect 31205 28611 31263 28617
rect 31205 28577 31217 28611
rect 31251 28608 31263 28611
rect 31754 28608 31760 28620
rect 31251 28580 31760 28608
rect 31251 28577 31263 28580
rect 31205 28571 31263 28577
rect 31754 28568 31760 28580
rect 31812 28608 31818 28620
rect 33042 28608 33048 28620
rect 31812 28580 33048 28608
rect 31812 28568 31818 28580
rect 33042 28568 33048 28580
rect 33100 28568 33106 28620
rect 40402 28568 40408 28620
rect 40460 28608 40466 28620
rect 40957 28611 41015 28617
rect 40957 28608 40969 28611
rect 40460 28580 40969 28608
rect 40460 28568 40466 28580
rect 40957 28577 40969 28580
rect 41003 28577 41015 28611
rect 40957 28571 41015 28577
rect 24765 28543 24823 28549
rect 24765 28509 24777 28543
rect 24811 28509 24823 28543
rect 25498 28540 25504 28552
rect 25459 28512 25504 28540
rect 24765 28503 24823 28509
rect 24780 28472 24808 28503
rect 25498 28500 25504 28512
rect 25556 28500 25562 28552
rect 26329 28543 26387 28549
rect 26329 28540 26341 28543
rect 26206 28512 26341 28540
rect 24946 28472 24952 28484
rect 24780 28444 24952 28472
rect 24946 28432 24952 28444
rect 25004 28472 25010 28484
rect 26206 28472 26234 28512
rect 26329 28509 26341 28512
rect 26375 28540 26387 28543
rect 29638 28540 29644 28552
rect 26375 28512 29644 28540
rect 26375 28509 26387 28512
rect 26329 28503 26387 28509
rect 29638 28500 29644 28512
rect 29696 28540 29702 28552
rect 29733 28543 29791 28549
rect 29733 28540 29745 28543
rect 29696 28512 29745 28540
rect 29696 28500 29702 28512
rect 29733 28509 29745 28512
rect 29779 28509 29791 28543
rect 29733 28503 29791 28509
rect 31389 28543 31447 28549
rect 31389 28509 31401 28543
rect 31435 28540 31447 28543
rect 31846 28540 31852 28552
rect 31435 28512 31852 28540
rect 31435 28509 31447 28512
rect 31389 28503 31447 28509
rect 31846 28500 31852 28512
rect 31904 28500 31910 28552
rect 35158 28540 35164 28552
rect 35119 28512 35164 28540
rect 35158 28500 35164 28512
rect 35216 28500 35222 28552
rect 35428 28543 35486 28549
rect 35428 28509 35440 28543
rect 35474 28540 35486 28543
rect 35894 28540 35900 28552
rect 35474 28512 35900 28540
rect 35474 28509 35486 28512
rect 35428 28503 35486 28509
rect 35894 28500 35900 28512
rect 35952 28500 35958 28552
rect 37001 28543 37059 28549
rect 37001 28509 37013 28543
rect 37047 28540 37059 28543
rect 40420 28540 40448 28568
rect 37047 28512 40448 28540
rect 40972 28540 41000 28571
rect 42797 28543 42855 28549
rect 42797 28540 42809 28543
rect 40972 28512 42809 28540
rect 37047 28509 37059 28512
rect 37001 28503 37059 28509
rect 42797 28509 42809 28512
rect 42843 28509 42855 28543
rect 42797 28503 42855 28509
rect 42886 28500 42892 28552
rect 42944 28540 42950 28552
rect 43053 28543 43111 28549
rect 43053 28540 43065 28543
rect 42944 28512 43065 28540
rect 42944 28500 42950 28512
rect 43053 28509 43065 28512
rect 43099 28509 43111 28543
rect 43053 28503 43111 28509
rect 25004 28444 26234 28472
rect 37268 28475 37326 28481
rect 25004 28432 25010 28444
rect 37268 28441 37280 28475
rect 37314 28472 37326 28475
rect 37918 28472 37924 28484
rect 37314 28444 37924 28472
rect 37314 28441 37326 28444
rect 37268 28435 37326 28441
rect 37918 28432 37924 28444
rect 37976 28432 37982 28484
rect 40862 28432 40868 28484
rect 40920 28472 40926 28484
rect 41202 28475 41260 28481
rect 41202 28472 41214 28475
rect 40920 28444 41214 28472
rect 40920 28432 40926 28444
rect 41202 28441 41214 28444
rect 41248 28441 41260 28475
rect 41202 28435 41260 28441
rect 26326 28404 26332 28416
rect 26287 28376 26332 28404
rect 26326 28364 26332 28376
rect 26384 28364 26390 28416
rect 29917 28407 29975 28413
rect 29917 28373 29929 28407
rect 29963 28404 29975 28407
rect 30190 28404 30196 28416
rect 29963 28376 30196 28404
rect 29963 28373 29975 28376
rect 29917 28367 29975 28373
rect 30190 28364 30196 28376
rect 30248 28364 30254 28416
rect 31386 28364 31392 28416
rect 31444 28404 31450 28416
rect 31573 28407 31631 28413
rect 31573 28404 31585 28407
rect 31444 28376 31585 28404
rect 31444 28364 31450 28376
rect 31573 28373 31585 28376
rect 31619 28373 31631 28407
rect 31573 28367 31631 28373
rect 31662 28364 31668 28416
rect 31720 28404 31726 28416
rect 38194 28404 38200 28416
rect 31720 28376 38200 28404
rect 31720 28364 31726 28376
rect 38194 28364 38200 28376
rect 38252 28404 38258 28416
rect 38381 28407 38439 28413
rect 38381 28404 38393 28407
rect 38252 28376 38393 28404
rect 38252 28364 38258 28376
rect 38381 28373 38393 28376
rect 38427 28373 38439 28407
rect 38381 28367 38439 28373
rect 41046 28364 41052 28416
rect 41104 28404 41110 28416
rect 42337 28407 42395 28413
rect 42337 28404 42349 28407
rect 41104 28376 42349 28404
rect 41104 28364 41110 28376
rect 42337 28373 42349 28376
rect 42383 28373 42395 28407
rect 42337 28367 42395 28373
rect 1104 28314 68816 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 68816 28314
rect 1104 28240 68816 28262
rect 31662 28200 31668 28212
rect 23032 28172 31668 28200
rect 23032 28073 23060 28172
rect 31662 28160 31668 28172
rect 31720 28160 31726 28212
rect 35158 28160 35164 28212
rect 35216 28200 35222 28212
rect 35529 28203 35587 28209
rect 35529 28200 35541 28203
rect 35216 28172 35541 28200
rect 35216 28160 35222 28172
rect 35529 28169 35541 28172
rect 35575 28169 35587 28203
rect 40862 28200 40868 28212
rect 40823 28172 40868 28200
rect 35529 28163 35587 28169
rect 40862 28160 40868 28172
rect 40920 28160 40926 28212
rect 25498 28092 25504 28144
rect 25556 28092 25562 28144
rect 27614 28092 27620 28144
rect 27672 28132 27678 28144
rect 27985 28135 28043 28141
rect 27985 28132 27997 28135
rect 27672 28104 27997 28132
rect 27672 28092 27678 28104
rect 27985 28101 27997 28104
rect 28031 28101 28043 28135
rect 27985 28095 28043 28101
rect 28201 28135 28259 28141
rect 28201 28101 28213 28135
rect 28247 28132 28259 28135
rect 28810 28132 28816 28144
rect 28247 28104 28672 28132
rect 28771 28104 28816 28132
rect 28247 28101 28259 28104
rect 28201 28095 28259 28101
rect 23017 28067 23075 28073
rect 23017 28033 23029 28067
rect 23063 28033 23075 28067
rect 25516 28064 25544 28092
rect 25685 28067 25743 28073
rect 25685 28064 25697 28067
rect 25516 28036 25697 28064
rect 23017 28027 23075 28033
rect 25685 28033 25697 28036
rect 25731 28033 25743 28067
rect 25685 28027 25743 28033
rect 25869 28067 25927 28073
rect 25869 28033 25881 28067
rect 25915 28064 25927 28067
rect 27157 28067 27215 28073
rect 27157 28064 27169 28067
rect 25915 28036 27169 28064
rect 25915 28033 25927 28036
rect 25869 28027 25927 28033
rect 27157 28033 27169 28036
rect 27203 28033 27215 28067
rect 28644 28064 28672 28104
rect 28810 28092 28816 28104
rect 28868 28092 28874 28144
rect 29029 28135 29087 28141
rect 29029 28132 29041 28135
rect 28920 28104 29041 28132
rect 28920 28064 28948 28104
rect 29029 28101 29041 28104
rect 29075 28132 29087 28135
rect 29730 28132 29736 28144
rect 29075 28104 29736 28132
rect 29075 28101 29087 28104
rect 29029 28095 29087 28101
rect 29730 28092 29736 28104
rect 29788 28092 29794 28144
rect 40402 28132 40408 28144
rect 38856 28104 40408 28132
rect 30190 28064 30196 28076
rect 28644 28036 28948 28064
rect 30151 28036 30196 28064
rect 27157 28027 27215 28033
rect 30190 28024 30196 28036
rect 30248 28024 30254 28076
rect 30460 28067 30518 28073
rect 30460 28033 30472 28067
rect 30506 28064 30518 28067
rect 31202 28064 31208 28076
rect 30506 28036 31208 28064
rect 30506 28033 30518 28036
rect 30460 28027 30518 28033
rect 31202 28024 31208 28036
rect 31260 28024 31266 28076
rect 33413 28067 33471 28073
rect 33413 28033 33425 28067
rect 33459 28064 33471 28067
rect 34790 28064 34796 28076
rect 33459 28036 34796 28064
rect 33459 28033 33471 28036
rect 33413 28027 33471 28033
rect 34790 28024 34796 28036
rect 34848 28024 34854 28076
rect 35345 28067 35403 28073
rect 35345 28033 35357 28067
rect 35391 28064 35403 28067
rect 35618 28064 35624 28076
rect 35391 28036 35624 28064
rect 35391 28033 35403 28036
rect 35345 28027 35403 28033
rect 23198 27996 23204 28008
rect 23159 27968 23204 27996
rect 23198 27956 23204 27968
rect 23256 27956 23262 28008
rect 23477 27999 23535 28005
rect 23477 27965 23489 27999
rect 23523 27965 23535 27999
rect 23477 27959 23535 27965
rect 25501 27999 25559 28005
rect 25501 27965 25513 27999
rect 25547 27996 25559 27999
rect 26510 27996 26516 28008
rect 25547 27968 26516 27996
rect 25547 27965 25559 27968
rect 25501 27959 25559 27965
rect 13814 27888 13820 27940
rect 13872 27928 13878 27940
rect 23492 27928 23520 27959
rect 26510 27956 26516 27968
rect 26568 27996 26574 28008
rect 27430 27996 27436 28008
rect 26568 27968 27436 27996
rect 26568 27956 26574 27968
rect 27430 27956 27436 27968
rect 27488 27956 27494 28008
rect 28902 27956 28908 28008
rect 28960 27996 28966 28008
rect 34057 27999 34115 28005
rect 34057 27996 34069 27999
rect 28960 27968 29316 27996
rect 28960 27956 28966 27968
rect 29086 27928 29092 27940
rect 13872 27900 23520 27928
rect 28184 27900 29092 27928
rect 13872 27888 13878 27900
rect 26602 27820 26608 27872
rect 26660 27860 26666 27872
rect 28184 27869 28212 27900
rect 26973 27863 27031 27869
rect 26973 27860 26985 27863
rect 26660 27832 26985 27860
rect 26660 27820 26666 27832
rect 26973 27829 26985 27832
rect 27019 27829 27031 27863
rect 26973 27823 27031 27829
rect 28169 27863 28227 27869
rect 28169 27829 28181 27863
rect 28215 27829 28227 27863
rect 28350 27860 28356 27872
rect 28311 27832 28356 27860
rect 28169 27823 28227 27829
rect 28350 27820 28356 27832
rect 28408 27820 28414 27872
rect 29012 27869 29040 27900
rect 29086 27888 29092 27900
rect 29144 27888 29150 27940
rect 28997 27863 29055 27869
rect 28997 27829 29009 27863
rect 29043 27829 29055 27863
rect 29178 27860 29184 27872
rect 29139 27832 29184 27860
rect 28997 27823 29055 27829
rect 29178 27820 29184 27832
rect 29236 27820 29242 27872
rect 29288 27860 29316 27968
rect 31211 27968 34069 27996
rect 31211 27860 31239 27968
rect 34057 27965 34069 27968
rect 34103 27965 34115 27999
rect 34330 27996 34336 28008
rect 34291 27968 34336 27996
rect 34057 27959 34115 27965
rect 34330 27956 34336 27968
rect 34388 27956 34394 28008
rect 34514 27956 34520 28008
rect 34572 27996 34578 28008
rect 35360 27996 35388 28027
rect 35618 28024 35624 28036
rect 35676 28024 35682 28076
rect 38856 28073 38884 28104
rect 40402 28092 40408 28104
rect 40460 28092 40466 28144
rect 44358 28132 44364 28144
rect 41248 28104 44364 28132
rect 39114 28073 39120 28076
rect 38841 28067 38899 28073
rect 38841 28033 38853 28067
rect 38887 28033 38899 28067
rect 39108 28064 39120 28073
rect 39075 28036 39120 28064
rect 38841 28027 38899 28033
rect 39108 28027 39120 28036
rect 39114 28024 39120 28027
rect 39172 28024 39178 28076
rect 40034 28024 40040 28076
rect 40092 28064 40098 28076
rect 41046 28064 41052 28076
rect 40092 28036 41052 28064
rect 40092 28024 40098 28036
rect 41046 28024 41052 28036
rect 41104 28064 41110 28076
rect 41248 28073 41276 28104
rect 44358 28092 44364 28104
rect 44416 28092 44422 28144
rect 41141 28067 41199 28073
rect 41141 28064 41153 28067
rect 41104 28036 41153 28064
rect 41104 28024 41110 28036
rect 41141 28033 41153 28036
rect 41187 28033 41199 28067
rect 41141 28027 41199 28033
rect 41233 28067 41291 28073
rect 41233 28033 41245 28067
rect 41279 28033 41291 28067
rect 41233 28027 41291 28033
rect 41325 28067 41383 28073
rect 41325 28033 41337 28067
rect 41371 28033 41383 28067
rect 41506 28064 41512 28076
rect 41467 28036 41512 28064
rect 41325 28027 41383 28033
rect 34572 27968 35388 27996
rect 34572 27956 34578 27968
rect 40678 27956 40684 28008
rect 40736 27996 40742 28008
rect 41340 27996 41368 28027
rect 41506 28024 41512 28036
rect 41564 28024 41570 28076
rect 40736 27968 41368 27996
rect 40736 27956 40742 27968
rect 31573 27931 31631 27937
rect 31573 27897 31585 27931
rect 31619 27928 31631 27931
rect 31754 27928 31760 27940
rect 31619 27900 31760 27928
rect 31619 27897 31631 27900
rect 31573 27891 31631 27897
rect 31754 27888 31760 27900
rect 31812 27888 31818 27940
rect 33226 27860 33232 27872
rect 29288 27832 31239 27860
rect 33187 27832 33232 27860
rect 33226 27820 33232 27832
rect 33284 27820 33290 27872
rect 40218 27860 40224 27872
rect 40179 27832 40224 27860
rect 40218 27820 40224 27832
rect 40276 27820 40282 27872
rect 1104 27770 68816 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 68816 27770
rect 1104 27696 68816 27718
rect 23198 27656 23204 27668
rect 23159 27628 23204 27656
rect 23198 27616 23204 27628
rect 23256 27616 23262 27668
rect 27614 27616 27620 27668
rect 27672 27656 27678 27668
rect 28353 27659 28411 27665
rect 28353 27656 28365 27659
rect 27672 27628 28365 27656
rect 27672 27616 27678 27628
rect 28353 27625 28365 27628
rect 28399 27625 28411 27659
rect 31202 27656 31208 27668
rect 31163 27628 31208 27656
rect 28353 27619 28411 27625
rect 31202 27616 31208 27628
rect 31260 27616 31266 27668
rect 38396 27628 38608 27656
rect 34054 27588 34060 27600
rect 34015 27560 34060 27588
rect 34054 27548 34060 27560
rect 34112 27588 34118 27600
rect 34112 27560 34744 27588
rect 34112 27548 34118 27560
rect 26142 27520 26148 27532
rect 26103 27492 26148 27520
rect 26142 27480 26148 27492
rect 26200 27480 26206 27532
rect 28810 27480 28816 27532
rect 28868 27520 28874 27532
rect 30006 27520 30012 27532
rect 28868 27492 30012 27520
rect 28868 27480 28874 27492
rect 30006 27480 30012 27492
rect 30064 27480 30070 27532
rect 34514 27520 34520 27532
rect 33888 27492 34520 27520
rect 23109 27455 23167 27461
rect 23109 27421 23121 27455
rect 23155 27452 23167 27455
rect 24302 27452 24308 27464
rect 23155 27424 24308 27452
rect 23155 27421 23167 27424
rect 23109 27415 23167 27421
rect 24302 27412 24308 27424
rect 24360 27412 24366 27464
rect 24397 27455 24455 27461
rect 24397 27421 24409 27455
rect 24443 27421 24455 27455
rect 26970 27452 26976 27464
rect 26931 27424 26976 27452
rect 24397 27415 24455 27421
rect 24412 27316 24440 27415
rect 26970 27412 26976 27424
rect 27028 27412 27034 27464
rect 28997 27455 29055 27461
rect 28997 27421 29009 27455
rect 29043 27452 29055 27455
rect 29178 27452 29184 27464
rect 29043 27424 29184 27452
rect 29043 27421 29055 27424
rect 28997 27415 29055 27421
rect 29178 27412 29184 27424
rect 29236 27412 29242 27464
rect 29733 27455 29791 27461
rect 29733 27421 29745 27455
rect 29779 27421 29791 27455
rect 30466 27452 30472 27464
rect 30427 27424 30472 27452
rect 29733 27415 29791 27421
rect 24578 27384 24584 27396
rect 24539 27356 24584 27384
rect 24578 27344 24584 27356
rect 24636 27344 24642 27396
rect 27240 27387 27298 27393
rect 27240 27353 27252 27387
rect 27286 27384 27298 27387
rect 27522 27384 27528 27396
rect 27286 27356 27528 27384
rect 27286 27353 27298 27356
rect 27240 27347 27298 27353
rect 27522 27344 27528 27356
rect 27580 27344 27586 27396
rect 27614 27344 27620 27396
rect 27672 27384 27678 27396
rect 29748 27384 29776 27415
rect 30466 27412 30472 27424
rect 30524 27412 30530 27464
rect 31386 27452 31392 27464
rect 31347 27424 31392 27452
rect 31386 27412 31392 27424
rect 31444 27412 31450 27464
rect 32674 27452 32680 27464
rect 32635 27424 32680 27452
rect 32674 27412 32680 27424
rect 32732 27412 32738 27464
rect 32944 27455 33002 27461
rect 32944 27421 32956 27455
rect 32990 27452 33002 27455
rect 33226 27452 33232 27464
rect 32990 27424 33232 27452
rect 32990 27421 33002 27424
rect 32944 27415 33002 27421
rect 33226 27412 33232 27424
rect 33284 27412 33290 27464
rect 33888 27384 33916 27492
rect 34514 27480 34520 27492
rect 34572 27480 34578 27532
rect 34716 27529 34744 27560
rect 34790 27548 34796 27600
rect 34848 27588 34854 27600
rect 35069 27591 35127 27597
rect 35069 27588 35081 27591
rect 34848 27560 35081 27588
rect 34848 27548 34854 27560
rect 35069 27557 35081 27560
rect 35115 27557 35127 27591
rect 38396 27588 38424 27628
rect 35069 27551 35127 27557
rect 37108 27560 38424 27588
rect 34701 27523 34759 27529
rect 34701 27489 34713 27523
rect 34747 27489 34759 27523
rect 34701 27483 34759 27489
rect 33962 27412 33968 27464
rect 34020 27452 34026 27464
rect 34330 27452 34336 27464
rect 34020 27424 34336 27452
rect 34020 27412 34026 27424
rect 34330 27412 34336 27424
rect 34388 27452 34394 27464
rect 34885 27455 34943 27461
rect 34885 27452 34897 27455
rect 34388 27424 34897 27452
rect 34388 27412 34394 27424
rect 34885 27421 34897 27424
rect 34931 27421 34943 27455
rect 34885 27415 34943 27421
rect 27672 27356 33916 27384
rect 27672 27344 27678 27356
rect 34238 27344 34244 27396
rect 34296 27384 34302 27396
rect 37108 27384 37136 27560
rect 38470 27548 38476 27600
rect 38528 27548 38534 27600
rect 38580 27588 38608 27628
rect 40218 27588 40224 27600
rect 38580 27560 40224 27588
rect 40218 27548 40224 27560
rect 40276 27548 40282 27600
rect 37185 27523 37243 27529
rect 37185 27489 37197 27523
rect 37231 27520 37243 27523
rect 38488 27520 38516 27548
rect 37231 27492 38516 27520
rect 38565 27523 38623 27529
rect 37231 27489 37243 27492
rect 37185 27483 37243 27489
rect 38565 27489 38577 27523
rect 38611 27489 38623 27523
rect 38565 27483 38623 27489
rect 37366 27384 37372 27396
rect 34296 27356 37136 27384
rect 37327 27356 37372 27384
rect 34296 27344 34302 27356
rect 37366 27344 37372 27356
rect 37424 27344 37430 27396
rect 28718 27316 28724 27328
rect 24412 27288 28724 27316
rect 28718 27276 28724 27288
rect 28776 27276 28782 27328
rect 28813 27319 28871 27325
rect 28813 27285 28825 27319
rect 28859 27316 28871 27319
rect 28902 27316 28908 27328
rect 28859 27288 28908 27316
rect 28859 27285 28871 27288
rect 28813 27279 28871 27285
rect 28902 27276 28908 27288
rect 28960 27276 28966 27328
rect 29730 27316 29736 27328
rect 29691 27288 29736 27316
rect 29730 27276 29736 27288
rect 29788 27276 29794 27328
rect 30650 27316 30656 27328
rect 30611 27288 30656 27316
rect 30650 27276 30656 27288
rect 30708 27276 30714 27328
rect 32858 27276 32864 27328
rect 32916 27316 32922 27328
rect 38580 27316 38608 27483
rect 40862 27452 40868 27464
rect 40823 27424 40868 27452
rect 40862 27412 40868 27424
rect 40920 27412 40926 27464
rect 32916 27288 38608 27316
rect 40957 27319 41015 27325
rect 32916 27276 32922 27288
rect 40957 27285 40969 27319
rect 41003 27316 41015 27319
rect 41506 27316 41512 27328
rect 41003 27288 41512 27316
rect 41003 27285 41015 27288
rect 40957 27279 41015 27285
rect 41506 27276 41512 27288
rect 41564 27276 41570 27328
rect 1104 27226 68816 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 68816 27226
rect 1104 27152 68816 27174
rect 24489 27115 24547 27121
rect 24489 27081 24501 27115
rect 24535 27112 24547 27115
rect 24578 27112 24584 27124
rect 24535 27084 24584 27112
rect 24535 27081 24547 27084
rect 24489 27075 24547 27081
rect 24578 27072 24584 27084
rect 24636 27072 24642 27124
rect 26421 27115 26479 27121
rect 26421 27081 26433 27115
rect 26467 27112 26479 27115
rect 26510 27112 26516 27124
rect 26467 27084 26516 27112
rect 26467 27081 26479 27084
rect 26421 27075 26479 27081
rect 26510 27072 26516 27084
rect 26568 27072 26574 27124
rect 26970 27072 26976 27124
rect 27028 27112 27034 27124
rect 27617 27115 27675 27121
rect 27617 27112 27629 27115
rect 27028 27084 27629 27112
rect 27028 27072 27034 27084
rect 27617 27081 27629 27084
rect 27663 27081 27675 27115
rect 27617 27075 27675 27081
rect 28718 27072 28724 27124
rect 28776 27112 28782 27124
rect 30006 27112 30012 27124
rect 28776 27084 29868 27112
rect 29967 27084 30012 27112
rect 28776 27072 28782 27084
rect 25308 27047 25366 27053
rect 25308 27013 25320 27047
rect 25354 27044 25366 27047
rect 26602 27044 26608 27056
rect 25354 27016 26608 27044
rect 25354 27013 25366 27016
rect 25308 27007 25366 27013
rect 26602 27004 26608 27016
rect 26660 27004 26666 27056
rect 29730 27044 29736 27056
rect 28644 27016 29736 27044
rect 24302 26936 24308 26988
rect 24360 26976 24366 26988
rect 24397 26979 24455 26985
rect 24397 26976 24409 26979
rect 24360 26948 24409 26976
rect 24360 26936 24366 26948
rect 24397 26945 24409 26948
rect 24443 26945 24455 26979
rect 24397 26939 24455 26945
rect 25041 26979 25099 26985
rect 25041 26945 25053 26979
rect 25087 26976 25099 26979
rect 26326 26976 26332 26988
rect 25087 26948 26332 26976
rect 25087 26945 25099 26948
rect 25041 26939 25099 26945
rect 26326 26936 26332 26948
rect 26384 26936 26390 26988
rect 27525 26979 27583 26985
rect 27525 26945 27537 26979
rect 27571 26976 27583 26979
rect 27614 26976 27620 26988
rect 27571 26948 27620 26976
rect 27571 26945 27583 26948
rect 27525 26939 27583 26945
rect 27614 26936 27620 26948
rect 27672 26936 27678 26988
rect 28644 26985 28672 27016
rect 29730 27004 29736 27016
rect 29788 27004 29794 27056
rect 29840 27044 29868 27084
rect 30006 27072 30012 27084
rect 30064 27072 30070 27124
rect 32674 27112 32680 27124
rect 32635 27084 32680 27112
rect 32674 27072 32680 27084
rect 32732 27072 32738 27124
rect 35526 27112 35532 27124
rect 34440 27084 35532 27112
rect 34238 27044 34244 27056
rect 29840 27016 34244 27044
rect 34238 27004 34244 27016
rect 34296 27004 34302 27056
rect 28902 26985 28908 26988
rect 28629 26979 28687 26985
rect 28629 26945 28641 26979
rect 28675 26945 28687 26979
rect 28896 26976 28908 26985
rect 28863 26948 28908 26976
rect 28629 26939 28687 26945
rect 28896 26939 28908 26948
rect 28902 26936 28908 26939
rect 28960 26936 28966 26988
rect 30650 26936 30656 26988
rect 30708 26976 30714 26988
rect 32493 26979 32551 26985
rect 32493 26976 32505 26979
rect 30708 26948 32505 26976
rect 30708 26936 30714 26948
rect 32493 26945 32505 26948
rect 32539 26945 32551 26979
rect 32493 26939 32551 26945
rect 33134 26936 33140 26988
rect 33192 26976 33198 26988
rect 33962 26976 33968 26988
rect 33192 26948 33968 26976
rect 33192 26936 33198 26948
rect 33962 26936 33968 26948
rect 34020 26936 34026 26988
rect 33781 26911 33839 26917
rect 33781 26877 33793 26911
rect 33827 26908 33839 26911
rect 34440 26908 34468 27084
rect 35526 27072 35532 27084
rect 35584 27112 35590 27124
rect 35989 27115 36047 27121
rect 35989 27112 36001 27115
rect 35584 27084 36001 27112
rect 35584 27072 35590 27084
rect 35989 27081 36001 27084
rect 36035 27081 36047 27115
rect 37366 27112 37372 27124
rect 37327 27084 37372 27112
rect 35989 27075 36047 27081
rect 37366 27072 37372 27084
rect 37424 27072 37430 27124
rect 33827 26880 34468 26908
rect 34532 27016 37320 27044
rect 33827 26877 33839 26880
rect 33781 26871 33839 26877
rect 34532 26840 34560 27016
rect 34609 26979 34667 26985
rect 34609 26945 34621 26979
rect 34655 26976 34667 26979
rect 34698 26976 34704 26988
rect 34655 26948 34704 26976
rect 34655 26945 34667 26948
rect 34609 26939 34667 26945
rect 34698 26936 34704 26948
rect 34756 26936 34762 26988
rect 34876 26979 34934 26985
rect 34876 26945 34888 26979
rect 34922 26976 34934 26979
rect 35434 26976 35440 26988
rect 34922 26948 35440 26976
rect 34922 26945 34934 26948
rect 34876 26939 34934 26945
rect 35434 26936 35440 26948
rect 35492 26936 35498 26988
rect 37292 26985 37320 27016
rect 37277 26979 37335 26985
rect 37277 26945 37289 26979
rect 37323 26945 37335 26979
rect 40034 26976 40040 26988
rect 39995 26948 40040 26976
rect 37277 26939 37335 26945
rect 31726 26812 34560 26840
rect 24210 26732 24216 26784
rect 24268 26772 24274 26784
rect 31726 26772 31754 26812
rect 24268 26744 31754 26772
rect 34149 26775 34207 26781
rect 24268 26732 24274 26744
rect 34149 26741 34161 26775
rect 34195 26772 34207 26775
rect 35618 26772 35624 26784
rect 34195 26744 35624 26772
rect 34195 26741 34207 26744
rect 34149 26735 34207 26741
rect 35618 26732 35624 26744
rect 35676 26732 35682 26784
rect 37292 26772 37320 26939
rect 40034 26936 40040 26948
rect 40092 26936 40098 26988
rect 40221 26911 40279 26917
rect 40221 26877 40233 26911
rect 40267 26908 40279 26911
rect 40310 26908 40316 26920
rect 40267 26880 40316 26908
rect 40267 26877 40279 26880
rect 40221 26871 40279 26877
rect 40310 26868 40316 26880
rect 40368 26868 40374 26920
rect 40497 26911 40555 26917
rect 40497 26877 40509 26911
rect 40543 26877 40555 26911
rect 40497 26871 40555 26877
rect 38838 26800 38844 26852
rect 38896 26840 38902 26852
rect 40512 26840 40540 26871
rect 38896 26812 40540 26840
rect 38896 26800 38902 26812
rect 45738 26772 45744 26784
rect 37292 26744 45744 26772
rect 45738 26732 45744 26744
rect 45796 26732 45802 26784
rect 1104 26682 68816 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 68816 26682
rect 1104 26608 68816 26630
rect 27522 26568 27528 26580
rect 27483 26540 27528 26568
rect 27522 26528 27528 26540
rect 27580 26528 27586 26580
rect 34698 26568 34704 26580
rect 31036 26540 34560 26568
rect 34659 26540 34704 26568
rect 24302 26460 24308 26512
rect 24360 26500 24366 26512
rect 31036 26500 31064 26540
rect 24360 26472 31064 26500
rect 32493 26503 32551 26509
rect 24360 26460 24366 26472
rect 32493 26469 32505 26503
rect 32539 26469 32551 26503
rect 32493 26463 32551 26469
rect 32508 26432 32536 26463
rect 32950 26432 32956 26444
rect 32508 26404 32956 26432
rect 32950 26392 32956 26404
rect 33008 26392 33014 26444
rect 34532 26432 34560 26540
rect 34698 26528 34704 26540
rect 34756 26528 34762 26580
rect 35434 26568 35440 26580
rect 35395 26540 35440 26568
rect 35434 26528 35440 26540
rect 35492 26528 35498 26580
rect 40310 26568 40316 26580
rect 40271 26540 40316 26568
rect 40310 26528 40316 26540
rect 40368 26528 40374 26580
rect 40862 26432 40868 26444
rect 34532 26404 40868 26432
rect 1670 26324 1676 26376
rect 1728 26364 1734 26376
rect 1949 26367 2007 26373
rect 1949 26364 1961 26367
rect 1728 26336 1961 26364
rect 1728 26324 1734 26336
rect 1949 26333 1961 26336
rect 1995 26333 2007 26367
rect 1949 26327 2007 26333
rect 3050 26324 3056 26376
rect 3108 26364 3114 26376
rect 27709 26367 27767 26373
rect 3108 26336 6914 26364
rect 3108 26324 3114 26336
rect 6886 26296 6914 26336
rect 27709 26333 27721 26367
rect 27755 26364 27767 26367
rect 28350 26364 28356 26376
rect 27755 26336 28356 26364
rect 27755 26333 27767 26336
rect 27709 26327 27767 26333
rect 28350 26324 28356 26336
rect 28408 26324 28414 26376
rect 31110 26364 31116 26376
rect 31071 26336 31116 26364
rect 31110 26324 31116 26336
rect 31168 26324 31174 26376
rect 32858 26364 32864 26376
rect 31211 26336 32864 26364
rect 31211 26296 31239 26336
rect 32858 26324 32864 26336
rect 32916 26324 32922 26376
rect 33134 26364 33140 26376
rect 33095 26336 33140 26364
rect 33134 26324 33140 26336
rect 33192 26324 33198 26376
rect 33778 26324 33784 26376
rect 33836 26364 33842 26376
rect 34701 26367 34759 26373
rect 34701 26364 34713 26367
rect 33836 26336 34713 26364
rect 33836 26324 33842 26336
rect 34701 26333 34713 26336
rect 34747 26333 34759 26367
rect 35618 26364 35624 26376
rect 35579 26336 35624 26364
rect 34701 26327 34759 26333
rect 35618 26324 35624 26336
rect 35676 26324 35682 26376
rect 40236 26373 40264 26404
rect 40862 26392 40868 26404
rect 40920 26392 40926 26444
rect 41230 26392 41236 26444
rect 41288 26432 41294 26444
rect 41325 26435 41383 26441
rect 41325 26432 41337 26435
rect 41288 26404 41337 26432
rect 41288 26392 41294 26404
rect 41325 26401 41337 26404
rect 41371 26401 41383 26435
rect 41506 26432 41512 26444
rect 41467 26404 41512 26432
rect 41325 26395 41383 26401
rect 41506 26392 41512 26404
rect 41564 26392 41570 26444
rect 40221 26367 40279 26373
rect 40221 26333 40233 26367
rect 40267 26333 40279 26367
rect 40221 26327 40279 26333
rect 6886 26268 31239 26296
rect 31380 26299 31438 26305
rect 31380 26265 31392 26299
rect 31426 26296 31438 26299
rect 32122 26296 32128 26308
rect 31426 26268 32128 26296
rect 31426 26265 31438 26268
rect 31380 26259 31438 26265
rect 32122 26256 32128 26268
rect 32180 26256 32186 26308
rect 43162 26296 43168 26308
rect 43123 26268 43168 26296
rect 43162 26256 43168 26268
rect 43220 26256 43226 26308
rect 33318 26228 33324 26240
rect 33279 26200 33324 26228
rect 33318 26188 33324 26200
rect 33376 26188 33382 26240
rect 1104 26138 68816 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 68816 26138
rect 1104 26064 68816 26086
rect 31110 26024 31116 26036
rect 31071 25996 31116 26024
rect 31110 25984 31116 25996
rect 31168 25984 31174 26036
rect 32122 26024 32128 26036
rect 32083 25996 32128 26024
rect 32122 25984 32128 25996
rect 32180 25984 32186 26036
rect 34790 25984 34796 26036
rect 34848 26024 34854 26036
rect 35069 26027 35127 26033
rect 35069 26024 35081 26027
rect 34848 25996 35081 26024
rect 34848 25984 34854 25996
rect 35069 25993 35081 25996
rect 35115 25993 35127 26027
rect 35069 25987 35127 25993
rect 30650 25916 30656 25968
rect 30708 25956 30714 25968
rect 31386 25956 31392 25968
rect 30708 25928 31392 25956
rect 30708 25916 30714 25928
rect 1670 25888 1676 25900
rect 1631 25860 1676 25888
rect 1670 25848 1676 25860
rect 1728 25848 1734 25900
rect 31128 25897 31156 25928
rect 31386 25916 31392 25928
rect 31444 25956 31450 25968
rect 33778 25956 33784 25968
rect 31444 25928 33784 25956
rect 31444 25916 31450 25928
rect 33778 25916 33784 25928
rect 33836 25916 33842 25968
rect 31113 25891 31171 25897
rect 31113 25857 31125 25891
rect 31159 25857 31171 25891
rect 31113 25851 31171 25857
rect 32309 25891 32367 25897
rect 32309 25857 32321 25891
rect 32355 25888 32367 25891
rect 33318 25888 33324 25900
rect 32355 25860 33324 25888
rect 32355 25857 32367 25860
rect 32309 25851 32367 25857
rect 33318 25848 33324 25860
rect 33376 25848 33382 25900
rect 33962 25897 33968 25900
rect 33956 25851 33968 25897
rect 34020 25888 34026 25900
rect 34020 25860 34056 25888
rect 33962 25848 33968 25851
rect 34020 25848 34026 25860
rect 1857 25823 1915 25829
rect 1857 25789 1869 25823
rect 1903 25820 1915 25823
rect 2314 25820 2320 25832
rect 1903 25792 2320 25820
rect 1903 25789 1915 25792
rect 1857 25783 1915 25789
rect 2314 25780 2320 25792
rect 2372 25780 2378 25832
rect 2774 25820 2780 25832
rect 2735 25792 2780 25820
rect 2774 25780 2780 25792
rect 2832 25780 2838 25832
rect 33686 25820 33692 25832
rect 33647 25792 33692 25820
rect 33686 25780 33692 25792
rect 33744 25780 33750 25832
rect 1104 25594 68816 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 68816 25594
rect 1104 25520 68816 25542
rect 2314 25480 2320 25492
rect 2275 25452 2320 25480
rect 2314 25440 2320 25452
rect 2372 25440 2378 25492
rect 33686 25440 33692 25492
rect 33744 25480 33750 25492
rect 33781 25483 33839 25489
rect 33781 25480 33793 25483
rect 33744 25452 33793 25480
rect 33744 25440 33750 25452
rect 33781 25449 33793 25452
rect 33827 25449 33839 25483
rect 33781 25443 33839 25449
rect 32490 25344 32496 25356
rect 32451 25316 32496 25344
rect 32490 25304 32496 25316
rect 32548 25304 32554 25356
rect 33152 25316 34928 25344
rect 33152 25288 33180 25316
rect 2225 25279 2283 25285
rect 2225 25245 2237 25279
rect 2271 25276 2283 25279
rect 3418 25276 3424 25288
rect 2271 25248 3424 25276
rect 2271 25245 2283 25248
rect 2225 25239 2283 25245
rect 3418 25236 3424 25248
rect 3476 25236 3482 25288
rect 32677 25279 32735 25285
rect 32677 25245 32689 25279
rect 32723 25276 32735 25279
rect 33134 25276 33140 25288
rect 32723 25248 33140 25276
rect 32723 25245 32735 25248
rect 32677 25239 32735 25245
rect 33134 25236 33140 25248
rect 33192 25236 33198 25288
rect 33778 25276 33784 25288
rect 33739 25248 33784 25276
rect 33778 25236 33784 25248
rect 33836 25236 33842 25288
rect 34790 25276 34796 25288
rect 34751 25248 34796 25276
rect 34790 25236 34796 25248
rect 34848 25236 34854 25288
rect 34900 25285 34928 25316
rect 34885 25279 34943 25285
rect 34885 25245 34897 25279
rect 34931 25245 34943 25279
rect 34885 25239 34943 25245
rect 32398 25100 32404 25152
rect 32456 25140 32462 25152
rect 32861 25143 32919 25149
rect 32861 25140 32873 25143
rect 32456 25112 32873 25140
rect 32456 25100 32462 25112
rect 32861 25109 32873 25112
rect 32907 25109 32919 25143
rect 35066 25140 35072 25152
rect 35027 25112 35072 25140
rect 32861 25103 32919 25109
rect 35066 25100 35072 25112
rect 35124 25100 35130 25152
rect 1104 25050 68816 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 68816 25050
rect 1104 24976 68816 24998
rect 33962 24896 33968 24948
rect 34020 24936 34026 24948
rect 34057 24939 34115 24945
rect 34057 24936 34069 24939
rect 34020 24908 34069 24936
rect 34020 24896 34026 24908
rect 34057 24905 34069 24908
rect 34103 24905 34115 24939
rect 34057 24899 34115 24905
rect 1854 24800 1860 24812
rect 1815 24772 1860 24800
rect 1854 24760 1860 24772
rect 1912 24760 1918 24812
rect 2593 24803 2651 24809
rect 2593 24769 2605 24803
rect 2639 24800 2651 24803
rect 5258 24800 5264 24812
rect 2639 24772 5264 24800
rect 2639 24769 2651 24772
rect 2593 24763 2651 24769
rect 5258 24760 5264 24772
rect 5316 24760 5322 24812
rect 31386 24800 31392 24812
rect 31347 24772 31392 24800
rect 31386 24760 31392 24772
rect 31444 24760 31450 24812
rect 32214 24760 32220 24812
rect 32272 24800 32278 24812
rect 32381 24803 32439 24809
rect 32381 24800 32393 24803
rect 32272 24772 32393 24800
rect 32272 24760 32278 24772
rect 32381 24769 32393 24772
rect 32427 24769 32439 24803
rect 32381 24763 32439 24769
rect 34241 24803 34299 24809
rect 34241 24769 34253 24803
rect 34287 24800 34299 24803
rect 35066 24800 35072 24812
rect 34287 24772 35072 24800
rect 34287 24769 34299 24772
rect 34241 24763 34299 24769
rect 35066 24760 35072 24772
rect 35124 24760 35130 24812
rect 2041 24735 2099 24741
rect 2041 24701 2053 24735
rect 2087 24732 2099 24735
rect 31481 24735 31539 24741
rect 2087 24704 6914 24732
rect 2087 24701 2099 24704
rect 2041 24695 2099 24701
rect 2038 24556 2044 24608
rect 2096 24596 2102 24608
rect 2685 24599 2743 24605
rect 2685 24596 2697 24599
rect 2096 24568 2697 24596
rect 2096 24556 2102 24568
rect 2685 24565 2697 24568
rect 2731 24565 2743 24599
rect 3418 24596 3424 24608
rect 3379 24568 3424 24596
rect 2685 24559 2743 24565
rect 3418 24556 3424 24568
rect 3476 24556 3482 24608
rect 6886 24596 6914 24704
rect 31481 24701 31493 24735
rect 31527 24732 31539 24735
rect 32125 24735 32183 24741
rect 32125 24732 32137 24735
rect 31527 24704 32137 24732
rect 31527 24701 31539 24704
rect 31481 24695 31539 24701
rect 32125 24701 32137 24704
rect 32171 24701 32183 24735
rect 32125 24695 32183 24701
rect 20714 24596 20720 24608
rect 6886 24568 20720 24596
rect 20714 24556 20720 24568
rect 20772 24556 20778 24608
rect 32490 24556 32496 24608
rect 32548 24596 32554 24608
rect 33505 24599 33563 24605
rect 33505 24596 33517 24599
rect 32548 24568 33517 24596
rect 32548 24556 32554 24568
rect 33505 24565 33517 24568
rect 33551 24565 33563 24599
rect 33505 24559 33563 24565
rect 1104 24506 68816 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 68816 24506
rect 1104 24432 68816 24454
rect 32214 24392 32220 24404
rect 32175 24364 32220 24392
rect 32214 24352 32220 24364
rect 32272 24352 32278 24404
rect 3418 24324 3424 24336
rect 1412 24296 3424 24324
rect 1412 24265 1440 24296
rect 3418 24284 3424 24296
rect 3476 24284 3482 24336
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24225 1455 24259
rect 1397 24219 1455 24225
rect 1581 24259 1639 24265
rect 1581 24225 1593 24259
rect 1627 24256 1639 24259
rect 2038 24256 2044 24268
rect 1627 24228 2044 24256
rect 1627 24225 1639 24228
rect 1581 24219 1639 24225
rect 2038 24216 2044 24228
rect 2096 24216 2102 24268
rect 2774 24256 2780 24268
rect 2735 24228 2780 24256
rect 2774 24216 2780 24228
rect 2832 24216 2838 24268
rect 32398 24188 32404 24200
rect 32359 24160 32404 24188
rect 32398 24148 32404 24160
rect 32456 24148 32462 24200
rect 1104 23962 68816 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 68816 23962
rect 1104 23888 68816 23910
rect 66254 23468 66260 23520
rect 66312 23508 66318 23520
rect 67637 23511 67695 23517
rect 67637 23508 67649 23511
rect 66312 23480 67649 23508
rect 66312 23468 66318 23480
rect 67637 23477 67649 23480
rect 67683 23477 67695 23511
rect 67637 23471 67695 23477
rect 1104 23418 68816 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 68816 23418
rect 1104 23344 68816 23366
rect 66254 23168 66260 23180
rect 66215 23140 66260 23168
rect 66254 23128 66260 23140
rect 66312 23128 66318 23180
rect 68094 23168 68100 23180
rect 68055 23140 68100 23168
rect 68094 23128 68100 23140
rect 68152 23128 68158 23180
rect 66438 23032 66444 23044
rect 66399 23004 66444 23032
rect 66438 22992 66444 23004
rect 66496 22992 66502 23044
rect 1104 22874 68816 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 68816 22874
rect 1104 22800 68816 22822
rect 66438 22720 66444 22772
rect 66496 22760 66502 22772
rect 67269 22763 67327 22769
rect 67269 22760 67281 22763
rect 66496 22732 67281 22760
rect 66496 22720 66502 22732
rect 67269 22729 67281 22732
rect 67315 22729 67327 22763
rect 67269 22723 67327 22729
rect 67174 22624 67180 22636
rect 67135 22596 67180 22624
rect 67174 22584 67180 22596
rect 67232 22584 67238 22636
rect 1762 22556 1768 22568
rect 1723 22528 1768 22556
rect 1762 22516 1768 22528
rect 1820 22516 1826 22568
rect 1949 22559 2007 22565
rect 1949 22525 1961 22559
rect 1995 22556 2007 22559
rect 2590 22556 2596 22568
rect 1995 22528 2596 22556
rect 1995 22525 2007 22528
rect 1949 22519 2007 22525
rect 2590 22516 2596 22528
rect 2648 22516 2654 22568
rect 2774 22556 2780 22568
rect 2735 22528 2780 22556
rect 2774 22516 2780 22528
rect 2832 22516 2838 22568
rect 1104 22330 68816 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 68816 22330
rect 1104 22256 68816 22278
rect 1762 22176 1768 22228
rect 1820 22216 1826 22228
rect 2041 22219 2099 22225
rect 2041 22216 2053 22219
rect 1820 22188 2053 22216
rect 1820 22176 1826 22188
rect 2041 22185 2053 22188
rect 2087 22185 2099 22219
rect 2590 22216 2596 22228
rect 2551 22188 2596 22216
rect 2041 22179 2099 22185
rect 2590 22176 2596 22188
rect 2648 22176 2654 22228
rect 66254 22108 66260 22160
rect 66312 22148 66318 22160
rect 67913 22151 67971 22157
rect 67913 22148 67925 22151
rect 66312 22120 67925 22148
rect 66312 22108 66318 22120
rect 67913 22117 67925 22120
rect 67959 22117 67971 22151
rect 67913 22111 67971 22117
rect 2501 22015 2559 22021
rect 2501 21981 2513 22015
rect 2547 22012 2559 22015
rect 4614 22012 4620 22024
rect 2547 21984 4620 22012
rect 2547 21981 2559 21984
rect 2501 21975 2559 21981
rect 4614 21972 4620 21984
rect 4672 21972 4678 22024
rect 1104 21786 68816 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 68816 21786
rect 1104 21712 68816 21734
rect 65978 21604 65984 21616
rect 65939 21576 65984 21604
rect 65978 21564 65984 21576
rect 66036 21564 66042 21616
rect 1854 21536 1860 21548
rect 1815 21508 1860 21536
rect 1854 21496 1860 21508
rect 1912 21496 1918 21548
rect 65797 21471 65855 21477
rect 65797 21437 65809 21471
rect 65843 21468 65855 21471
rect 66254 21468 66260 21480
rect 65843 21440 66260 21468
rect 65843 21437 65855 21440
rect 65797 21431 65855 21437
rect 66254 21428 66260 21440
rect 66312 21428 66318 21480
rect 67542 21468 67548 21480
rect 67503 21440 67548 21468
rect 67542 21428 67548 21440
rect 67600 21428 67606 21480
rect 1949 21335 2007 21341
rect 1949 21301 1961 21335
rect 1995 21332 2007 21335
rect 19150 21332 19156 21344
rect 1995 21304 19156 21332
rect 1995 21301 2007 21304
rect 1949 21295 2007 21301
rect 19150 21292 19156 21304
rect 19208 21292 19214 21344
rect 1104 21242 68816 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 68816 21242
rect 1104 21168 68816 21190
rect 1104 20698 68816 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 68816 20698
rect 1104 20624 68816 20646
rect 1104 20154 68816 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 68816 20154
rect 1104 20080 68816 20102
rect 1104 19610 68816 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 68816 19610
rect 1104 19536 68816 19558
rect 1104 19066 68816 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 68816 19066
rect 1104 18992 68816 19014
rect 67818 18748 67824 18760
rect 67779 18720 67824 18748
rect 67818 18708 67824 18720
rect 67876 18708 67882 18760
rect 68002 18612 68008 18624
rect 67963 18584 68008 18612
rect 68002 18572 68008 18584
rect 68060 18572 68066 18624
rect 1104 18522 68816 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 68816 18522
rect 1104 18448 68816 18470
rect 27709 18343 27767 18349
rect 27709 18309 27721 18343
rect 27755 18340 27767 18343
rect 28718 18340 28724 18352
rect 27755 18312 28724 18340
rect 27755 18309 27767 18312
rect 27709 18303 27767 18309
rect 28718 18300 28724 18312
rect 28776 18300 28782 18352
rect 26973 18275 27031 18281
rect 26973 18241 26985 18275
rect 27019 18272 27031 18275
rect 68002 18272 68008 18284
rect 27019 18244 68008 18272
rect 27019 18241 27031 18244
rect 26973 18235 27031 18241
rect 68002 18232 68008 18244
rect 68060 18232 68066 18284
rect 27341 18207 27399 18213
rect 27341 18173 27353 18207
rect 27387 18204 27399 18207
rect 27430 18204 27436 18216
rect 27387 18176 27436 18204
rect 27387 18173 27399 18176
rect 27341 18167 27399 18173
rect 27430 18164 27436 18176
rect 27488 18164 27494 18216
rect 3970 18096 3976 18148
rect 4028 18136 4034 18148
rect 27249 18139 27307 18145
rect 27249 18136 27261 18139
rect 4028 18108 27261 18136
rect 4028 18096 4034 18108
rect 27249 18105 27261 18108
rect 27295 18105 27307 18139
rect 27249 18099 27307 18105
rect 27138 18071 27196 18077
rect 27138 18037 27150 18071
rect 27184 18068 27196 18071
rect 36906 18068 36912 18080
rect 27184 18040 36912 18068
rect 27184 18037 27196 18040
rect 27138 18031 27196 18037
rect 36906 18028 36912 18040
rect 36964 18028 36970 18080
rect 1104 17978 68816 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 68816 17978
rect 1104 17904 68816 17926
rect 65794 17620 65800 17672
rect 65852 17660 65858 17672
rect 67913 17663 67971 17669
rect 67913 17660 67925 17663
rect 65852 17632 67925 17660
rect 65852 17620 65858 17632
rect 67913 17629 67925 17632
rect 67959 17629 67971 17663
rect 67913 17623 67971 17629
rect 1104 17434 68816 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 68816 17434
rect 1104 17360 68816 17382
rect 65981 17255 66039 17261
rect 65981 17221 65993 17255
rect 66027 17252 66039 17255
rect 67726 17252 67732 17264
rect 66027 17224 67732 17252
rect 66027 17221 66039 17224
rect 65981 17215 66039 17221
rect 67726 17212 67732 17224
rect 67784 17212 67790 17264
rect 65794 17184 65800 17196
rect 65755 17156 65800 17184
rect 65794 17144 65800 17156
rect 65852 17144 65858 17196
rect 67542 17116 67548 17128
rect 67503 17088 67548 17116
rect 67542 17076 67548 17088
rect 67600 17076 67606 17128
rect 1104 16890 68816 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 68816 16890
rect 1104 16816 68816 16838
rect 66714 16600 66720 16652
rect 66772 16640 66778 16652
rect 66772 16612 67588 16640
rect 66772 16600 66778 16612
rect 43162 16532 43168 16584
rect 43220 16572 43226 16584
rect 66162 16572 66168 16584
rect 43220 16544 66168 16572
rect 43220 16532 43226 16544
rect 66162 16532 66168 16544
rect 66220 16532 66226 16584
rect 67560 16581 67588 16612
rect 67545 16575 67603 16581
rect 67545 16541 67557 16575
rect 67591 16574 67603 16575
rect 67591 16546 67625 16574
rect 67591 16541 67603 16546
rect 67545 16535 67603 16541
rect 67637 16439 67695 16445
rect 67637 16405 67649 16439
rect 67683 16436 67695 16439
rect 67726 16436 67732 16448
rect 67683 16408 67732 16436
rect 67683 16405 67695 16408
rect 67637 16399 67695 16405
rect 67726 16396 67732 16408
rect 67784 16396 67790 16448
rect 1104 16346 68816 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 68816 16346
rect 1104 16272 68816 16294
rect 2038 16028 2044 16040
rect 1999 16000 2044 16028
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 2225 16031 2283 16037
rect 2225 15997 2237 16031
rect 2271 16028 2283 16031
rect 2866 16028 2872 16040
rect 2271 16000 2872 16028
rect 2271 15997 2283 16000
rect 2225 15991 2283 15997
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 2958 15988 2964 16040
rect 3016 16028 3022 16040
rect 3016 16000 3061 16028
rect 3016 15988 3022 16000
rect 1104 15802 68816 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 68816 15802
rect 1104 15728 68816 15750
rect 2038 15648 2044 15700
rect 2096 15688 2102 15700
rect 2317 15691 2375 15697
rect 2317 15688 2329 15691
rect 2096 15660 2329 15688
rect 2096 15648 2102 15660
rect 2317 15657 2329 15660
rect 2363 15657 2375 15691
rect 2866 15688 2872 15700
rect 2827 15660 2872 15688
rect 2317 15651 2375 15657
rect 2866 15648 2872 15660
rect 2924 15648 2930 15700
rect 2777 15487 2835 15493
rect 2777 15453 2789 15487
rect 2823 15484 2835 15487
rect 2866 15484 2872 15496
rect 2823 15456 2872 15484
rect 2823 15453 2835 15456
rect 2777 15447 2835 15453
rect 2866 15444 2872 15456
rect 2924 15484 2930 15496
rect 4706 15484 4712 15496
rect 2924 15456 4712 15484
rect 2924 15444 2930 15456
rect 4706 15444 4712 15456
rect 4764 15444 4770 15496
rect 67266 15444 67272 15496
rect 67324 15484 67330 15496
rect 67545 15487 67603 15493
rect 67545 15484 67557 15487
rect 67324 15456 67557 15484
rect 67324 15444 67330 15456
rect 67545 15453 67557 15456
rect 67591 15453 67603 15487
rect 67545 15447 67603 15453
rect 66254 15308 66260 15360
rect 66312 15348 66318 15360
rect 67637 15351 67695 15357
rect 67637 15348 67649 15351
rect 66312 15320 67649 15348
rect 66312 15308 66318 15320
rect 67637 15317 67649 15320
rect 67683 15317 67695 15351
rect 67637 15311 67695 15317
rect 1104 15258 68816 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 68816 15258
rect 1104 15184 68816 15206
rect 65981 15079 66039 15085
rect 65981 15045 65993 15079
rect 66027 15076 66039 15079
rect 66254 15076 66260 15088
rect 66027 15048 66260 15076
rect 66027 15045 66039 15048
rect 65981 15039 66039 15045
rect 66254 15036 66260 15048
rect 66312 15036 66318 15088
rect 65797 14943 65855 14949
rect 65797 14909 65809 14943
rect 65843 14940 65855 14943
rect 67358 14940 67364 14952
rect 65843 14912 67364 14940
rect 65843 14909 65855 14912
rect 65797 14903 65855 14909
rect 67358 14900 67364 14912
rect 67416 14900 67422 14952
rect 67542 14940 67548 14952
rect 67503 14912 67548 14940
rect 67542 14900 67548 14912
rect 67600 14900 67606 14952
rect 1104 14714 68816 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 68816 14714
rect 1104 14640 68816 14662
rect 67358 14560 67364 14612
rect 67416 14600 67422 14612
rect 67913 14603 67971 14609
rect 67913 14600 67925 14603
rect 67416 14572 67925 14600
rect 67416 14560 67422 14572
rect 67913 14569 67925 14572
rect 67959 14569 67971 14603
rect 67913 14563 67971 14569
rect 1104 14170 68816 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 68816 14170
rect 1104 14096 68816 14118
rect 1104 13626 68816 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 68816 13626
rect 1104 13552 68816 13574
rect 1578 13268 1584 13320
rect 1636 13308 1642 13320
rect 1765 13311 1823 13317
rect 1765 13308 1777 13311
rect 1636 13280 1777 13308
rect 1636 13268 1642 13280
rect 1765 13277 1777 13280
rect 1811 13277 1823 13311
rect 67818 13308 67824 13320
rect 67779 13280 67824 13308
rect 1765 13271 1823 13277
rect 67818 13268 67824 13280
rect 67876 13268 67882 13320
rect 68002 13172 68008 13184
rect 67963 13144 68008 13172
rect 68002 13132 68008 13144
rect 68060 13132 68066 13184
rect 1104 13082 68816 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 68816 13082
rect 1104 13008 68816 13030
rect 1578 12832 1584 12844
rect 1539 12804 1584 12832
rect 1578 12792 1584 12804
rect 1636 12792 1642 12844
rect 32122 12832 32128 12844
rect 32083 12804 32128 12832
rect 32122 12792 32128 12804
rect 32180 12792 32186 12844
rect 33137 12835 33195 12841
rect 33137 12832 33149 12835
rect 32416 12804 33149 12832
rect 1762 12764 1768 12776
rect 1723 12736 1768 12764
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 2774 12764 2780 12776
rect 2735 12736 2780 12764
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 31938 12724 31944 12776
rect 31996 12764 32002 12776
rect 32272 12767 32330 12773
rect 32272 12764 32284 12767
rect 31996 12736 32284 12764
rect 31996 12724 32002 12736
rect 32272 12733 32284 12736
rect 32318 12764 32330 12767
rect 32416 12764 32444 12804
rect 33137 12801 33149 12804
rect 33183 12801 33195 12835
rect 33137 12795 33195 12801
rect 32318 12736 32444 12764
rect 32493 12767 32551 12773
rect 32318 12733 32330 12736
rect 32272 12727 32330 12733
rect 32493 12733 32505 12767
rect 32539 12764 32551 12767
rect 68002 12764 68008 12776
rect 32539 12736 68008 12764
rect 32539 12733 32551 12736
rect 32493 12727 32551 12733
rect 68002 12724 68008 12736
rect 68060 12724 68066 12776
rect 32585 12699 32643 12705
rect 32585 12696 32597 12699
rect 26206 12668 32597 12696
rect 22554 12588 22560 12640
rect 22612 12628 22618 12640
rect 26206 12628 26234 12668
rect 32585 12665 32597 12668
rect 32631 12665 32643 12699
rect 32585 12659 32643 12665
rect 22612 12600 26234 12628
rect 22612 12588 22618 12600
rect 32398 12588 32404 12640
rect 32456 12628 32462 12640
rect 32456 12600 32501 12628
rect 32456 12588 32462 12600
rect 1104 12538 68816 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 68816 12538
rect 1104 12464 68816 12486
rect 1762 12384 1768 12436
rect 1820 12424 1826 12436
rect 2133 12427 2191 12433
rect 2133 12424 2145 12427
rect 1820 12396 2145 12424
rect 1820 12384 1826 12396
rect 2133 12393 2145 12396
rect 2179 12393 2191 12427
rect 2133 12387 2191 12393
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12220 2099 12223
rect 2406 12220 2412 12232
rect 2087 12192 2412 12220
rect 2087 12189 2099 12192
rect 2041 12183 2099 12189
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 1104 11994 68816 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 68816 11994
rect 1104 11920 68816 11942
rect 1104 11450 68816 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 68816 11450
rect 1104 11376 68816 11398
rect 1104 10906 68816 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 68816 10906
rect 1104 10832 68816 10854
rect 1104 10362 68816 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 68816 10362
rect 1104 10288 68816 10310
rect 1104 9818 68816 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 68816 9818
rect 1104 9744 68816 9766
rect 1104 9274 68816 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 68816 9274
rect 1104 9200 68816 9222
rect 1104 8730 68816 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 68816 8730
rect 1104 8656 68816 8678
rect 1104 8186 68816 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 68816 8186
rect 1104 8112 68816 8134
rect 67634 7868 67640 7880
rect 67595 7840 67640 7868
rect 67634 7828 67640 7840
rect 67692 7828 67698 7880
rect 1854 7800 1860 7812
rect 1815 7772 1860 7800
rect 1854 7760 1860 7772
rect 1912 7760 1918 7812
rect 19978 7760 19984 7812
rect 20036 7800 20042 7812
rect 67913 7803 67971 7809
rect 67913 7800 67925 7803
rect 20036 7772 67925 7800
rect 20036 7760 20042 7772
rect 67913 7769 67925 7772
rect 67959 7769 67971 7803
rect 67913 7763 67971 7769
rect 2133 7735 2191 7741
rect 2133 7701 2145 7735
rect 2179 7732 2191 7735
rect 17586 7732 17592 7744
rect 2179 7704 17592 7732
rect 2179 7701 2191 7704
rect 2133 7695 2191 7701
rect 17586 7692 17592 7704
rect 17644 7692 17650 7744
rect 1104 7642 68816 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 68816 7642
rect 1104 7568 68816 7590
rect 1104 7098 68816 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 68816 7098
rect 1104 7024 68816 7046
rect 65794 6740 65800 6792
rect 65852 6780 65858 6792
rect 67913 6783 67971 6789
rect 67913 6780 67925 6783
rect 65852 6752 67925 6780
rect 65852 6740 65858 6752
rect 67913 6749 67925 6752
rect 67959 6749 67971 6783
rect 67913 6743 67971 6749
rect 1104 6554 68816 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 68816 6554
rect 1104 6480 68816 6502
rect 65794 6304 65800 6316
rect 65755 6276 65800 6304
rect 65794 6264 65800 6276
rect 65852 6264 65858 6316
rect 65978 6236 65984 6248
rect 65939 6208 65984 6236
rect 65978 6196 65984 6208
rect 66036 6196 66042 6248
rect 67542 6236 67548 6248
rect 67503 6208 67548 6236
rect 67542 6196 67548 6208
rect 67600 6196 67606 6248
rect 1104 6010 68816 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 68816 6010
rect 1104 5936 68816 5958
rect 65978 5856 65984 5908
rect 66036 5896 66042 5908
rect 67637 5899 67695 5905
rect 67637 5896 67649 5899
rect 66036 5868 67649 5896
rect 66036 5856 66042 5868
rect 67637 5865 67649 5868
rect 67683 5865 67695 5899
rect 67637 5859 67695 5865
rect 45526 5732 66944 5760
rect 2774 5652 2780 5704
rect 2832 5692 2838 5704
rect 45526 5692 45554 5732
rect 66438 5692 66444 5704
rect 2832 5664 45554 5692
rect 66399 5664 66444 5692
rect 2832 5652 2838 5664
rect 66438 5652 66444 5664
rect 66496 5652 66502 5704
rect 66916 5701 66944 5732
rect 66901 5695 66959 5701
rect 66901 5661 66913 5695
rect 66947 5692 66959 5695
rect 67266 5692 67272 5704
rect 66947 5664 67272 5692
rect 66947 5661 66959 5664
rect 66901 5655 66959 5661
rect 67266 5652 67272 5664
rect 67324 5692 67330 5704
rect 67545 5695 67603 5701
rect 67545 5692 67557 5695
rect 67324 5664 67557 5692
rect 67324 5652 67330 5664
rect 67545 5661 67557 5664
rect 67591 5661 67603 5695
rect 67545 5655 67603 5661
rect 66990 5556 66996 5568
rect 66951 5528 66996 5556
rect 66990 5516 66996 5528
rect 67048 5516 67054 5568
rect 1104 5466 68816 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 68816 5466
rect 1104 5392 68816 5414
rect 65981 5287 66039 5293
rect 65981 5253 65993 5287
rect 66027 5284 66039 5287
rect 66990 5284 66996 5296
rect 66027 5256 66996 5284
rect 66027 5253 66039 5256
rect 65981 5247 66039 5253
rect 66990 5244 66996 5256
rect 67048 5244 67054 5296
rect 65797 5151 65855 5157
rect 65797 5117 65809 5151
rect 65843 5148 65855 5151
rect 66438 5148 66444 5160
rect 65843 5120 66444 5148
rect 65843 5117 65855 5120
rect 65797 5111 65855 5117
rect 66438 5108 66444 5120
rect 66496 5108 66502 5160
rect 67542 5148 67548 5160
rect 67503 5120 67548 5148
rect 67542 5108 67548 5120
rect 67600 5108 67606 5160
rect 1104 4922 68816 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 68816 4922
rect 1104 4848 68816 4870
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4604 5687 4607
rect 24118 4604 24124 4616
rect 5675 4576 24124 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 24118 4564 24124 4576
rect 24176 4564 24182 4616
rect 66898 4604 66904 4616
rect 66859 4576 66904 4604
rect 66898 4564 66904 4576
rect 66956 4564 66962 4616
rect 67266 4564 67272 4616
rect 67324 4604 67330 4616
rect 67361 4607 67419 4613
rect 67361 4604 67373 4607
rect 67324 4576 67373 4604
rect 67324 4564 67330 4576
rect 67361 4573 67373 4576
rect 67407 4573 67419 4607
rect 67361 4567 67419 4573
rect 6362 4496 6368 4548
rect 6420 4536 6426 4548
rect 10226 4536 10232 4548
rect 6420 4508 10232 4536
rect 6420 4496 6426 4508
rect 10226 4496 10232 4508
rect 10284 4496 10290 4548
rect 67450 4468 67456 4480
rect 67411 4440 67456 4468
rect 67450 4428 67456 4440
rect 67508 4428 67514 4480
rect 1104 4378 68816 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 68816 4378
rect 1104 4304 68816 4326
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 6362 4128 6368 4140
rect 5123 4100 6368 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 6822 4128 6828 4140
rect 6783 4100 6828 4128
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 34606 4088 34612 4140
rect 34664 4128 34670 4140
rect 36078 4128 36084 4140
rect 34664 4100 36084 4128
rect 34664 4088 34670 4100
rect 36078 4088 36084 4100
rect 36136 4088 36142 4140
rect 45738 4128 45744 4140
rect 45699 4100 45744 4128
rect 45738 4088 45744 4100
rect 45796 4088 45802 4140
rect 61933 4131 61991 4137
rect 61933 4097 61945 4131
rect 61979 4128 61991 4131
rect 61979 4100 64874 4128
rect 61979 4097 61991 4100
rect 61933 4091 61991 4097
rect 41230 4020 41236 4072
rect 41288 4060 41294 4072
rect 45922 4060 45928 4072
rect 41288 4032 45928 4060
rect 41288 4020 41294 4032
rect 45922 4020 45928 4032
rect 45980 4020 45986 4072
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 1857 3927 1915 3933
rect 1857 3924 1869 3927
rect 1636 3896 1869 3924
rect 1636 3884 1642 3896
rect 1857 3893 1869 3896
rect 1903 3893 1915 3927
rect 4614 3924 4620 3936
rect 4575 3896 4620 3924
rect 1857 3887 1915 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 5166 3924 5172 3936
rect 5127 3896 5172 3924
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 6822 3884 6828 3936
rect 6880 3924 6886 3936
rect 6917 3927 6975 3933
rect 6917 3924 6929 3927
rect 6880 3896 6929 3924
rect 6880 3884 6886 3896
rect 6917 3893 6929 3896
rect 6963 3893 6975 3927
rect 6917 3887 6975 3893
rect 45833 3927 45891 3933
rect 45833 3893 45845 3927
rect 45879 3924 45891 3927
rect 46382 3924 46388 3936
rect 45879 3896 46388 3924
rect 45879 3893 45891 3896
rect 45833 3887 45891 3893
rect 46382 3884 46388 3896
rect 46440 3884 46446 3936
rect 60642 3884 60648 3936
rect 60700 3924 60706 3936
rect 60921 3927 60979 3933
rect 60921 3924 60933 3927
rect 60700 3896 60933 3924
rect 60700 3884 60706 3896
rect 60921 3893 60933 3896
rect 60967 3893 60979 3927
rect 60921 3887 60979 3893
rect 62025 3927 62083 3933
rect 62025 3893 62037 3927
rect 62071 3924 62083 3927
rect 62114 3924 62120 3936
rect 62071 3896 62120 3924
rect 62071 3893 62083 3896
rect 62025 3887 62083 3893
rect 62114 3884 62120 3896
rect 62172 3884 62178 3936
rect 64846 3924 64874 4100
rect 65797 4063 65855 4069
rect 65797 4029 65809 4063
rect 65843 4029 65855 4063
rect 65797 4023 65855 4029
rect 65981 4063 66039 4069
rect 65981 4029 65993 4063
rect 66027 4060 66039 4063
rect 67450 4060 67456 4072
rect 66027 4032 67456 4060
rect 66027 4029 66039 4032
rect 65981 4023 66039 4029
rect 65812 3992 65840 4023
rect 67450 4020 67456 4032
rect 67508 4020 67514 4072
rect 67637 4063 67695 4069
rect 67637 4029 67649 4063
rect 67683 4060 67695 4063
rect 68922 4060 68928 4072
rect 67683 4032 68928 4060
rect 67683 4029 67695 4032
rect 67637 4023 67695 4029
rect 68922 4020 68928 4032
rect 68980 4020 68986 4072
rect 66898 3992 66904 4004
rect 65812 3964 66904 3992
rect 66898 3952 66904 3964
rect 66956 3952 66962 4004
rect 67174 3924 67180 3936
rect 64846 3896 67180 3924
rect 67174 3884 67180 3896
rect 67232 3884 67238 3936
rect 1104 3834 68816 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 68816 3834
rect 1104 3760 68816 3782
rect 658 3680 664 3732
rect 716 3720 722 3732
rect 716 3692 6914 3720
rect 716 3680 722 3692
rect 3142 3612 3148 3664
rect 3200 3652 3206 3664
rect 6886 3652 6914 3692
rect 47670 3652 47676 3664
rect 3200 3624 4936 3652
rect 6886 3624 47676 3652
rect 3200 3612 3206 3624
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3584 4491 3587
rect 4614 3584 4620 3596
rect 4479 3556 4620 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 4908 3593 4936 3624
rect 47670 3612 47676 3624
rect 47728 3612 47734 3664
rect 4893 3587 4951 3593
rect 4893 3553 4905 3587
rect 4939 3553 4951 3587
rect 10962 3584 10968 3596
rect 4893 3547 4951 3553
rect 6886 3556 7696 3584
rect 10923 3556 10968 3584
rect 1946 3516 1952 3528
rect 1907 3488 1952 3516
rect 1946 3476 1952 3488
rect 2004 3476 2010 3528
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3516 2835 3519
rect 3878 3516 3884 3528
rect 2823 3488 3884 3516
rect 2823 3485 2835 3488
rect 2777 3479 2835 3485
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 6733 3519 6791 3525
rect 6733 3485 6745 3519
rect 6779 3516 6791 3519
rect 6886 3516 6914 3556
rect 6779 3488 6914 3516
rect 7561 3519 7619 3525
rect 6779 3485 6791 3488
rect 6733 3479 6791 3485
rect 7561 3485 7573 3519
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 4617 3451 4675 3457
rect 4617 3417 4629 3451
rect 4663 3448 4675 3451
rect 5166 3448 5172 3460
rect 4663 3420 5172 3448
rect 4663 3417 4675 3420
rect 4617 3411 4675 3417
rect 5166 3408 5172 3420
rect 5224 3408 5230 3460
rect 6638 3408 6644 3460
rect 6696 3448 6702 3460
rect 7576 3448 7604 3479
rect 6696 3420 7604 3448
rect 6696 3408 6702 3420
rect 1762 3340 1768 3392
rect 1820 3380 1826 3392
rect 2041 3383 2099 3389
rect 2041 3380 2053 3383
rect 1820 3352 2053 3380
rect 1820 3340 1826 3352
rect 2041 3349 2053 3352
rect 2087 3349 2099 3383
rect 2041 3343 2099 3349
rect 6546 3340 6552 3392
rect 6604 3380 6610 3392
rect 6825 3383 6883 3389
rect 6825 3380 6837 3383
rect 6604 3352 6837 3380
rect 6604 3340 6610 3352
rect 6825 3349 6837 3352
rect 6871 3349 6883 3383
rect 7668 3380 7696 3556
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 16546 3556 22048 3584
rect 10410 3516 10416 3528
rect 10371 3488 10416 3516
rect 10410 3476 10416 3488
rect 10468 3476 10474 3528
rect 10594 3448 10600 3460
rect 10555 3420 10600 3448
rect 10594 3408 10600 3420
rect 10652 3408 10658 3460
rect 16546 3380 16574 3556
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 22020 3525 22048 3556
rect 23106 3544 23112 3596
rect 23164 3584 23170 3596
rect 46382 3584 46388 3596
rect 23164 3556 45048 3584
rect 46343 3556 46388 3584
rect 23164 3544 23170 3556
rect 19613 3519 19671 3525
rect 19613 3516 19625 3519
rect 19392 3488 19625 3516
rect 19392 3476 19398 3488
rect 19613 3485 19625 3488
rect 19659 3485 19671 3519
rect 19613 3479 19671 3485
rect 22005 3519 22063 3525
rect 22005 3485 22017 3519
rect 22051 3516 22063 3519
rect 23842 3516 23848 3528
rect 22051 3488 23848 3516
rect 22051 3485 22063 3488
rect 22005 3479 22063 3485
rect 23842 3476 23848 3488
rect 23900 3476 23906 3528
rect 38102 3476 38108 3528
rect 38160 3516 38166 3528
rect 45020 3525 45048 3556
rect 46382 3544 46388 3556
rect 46440 3544 46446 3596
rect 47026 3584 47032 3596
rect 46987 3556 47032 3584
rect 47026 3544 47032 3556
rect 47084 3544 47090 3596
rect 62114 3584 62120 3596
rect 62075 3556 62120 3584
rect 62114 3544 62120 3556
rect 62172 3544 62178 3596
rect 62482 3584 62488 3596
rect 62443 3556 62488 3584
rect 62482 3544 62488 3556
rect 62540 3544 62546 3596
rect 38381 3519 38439 3525
rect 38381 3516 38393 3519
rect 38160 3488 38393 3516
rect 38160 3476 38166 3488
rect 38381 3485 38393 3488
rect 38427 3485 38439 3519
rect 38381 3479 38439 3485
rect 45005 3519 45063 3525
rect 45005 3485 45017 3519
rect 45051 3485 45063 3519
rect 46198 3516 46204 3528
rect 46159 3488 46204 3516
rect 45005 3479 45063 3485
rect 46198 3476 46204 3488
rect 46256 3476 46262 3528
rect 50890 3476 50896 3528
rect 50948 3516 50954 3528
rect 51718 3516 51724 3528
rect 50948 3488 51724 3516
rect 50948 3476 50954 3488
rect 51718 3476 51724 3488
rect 51776 3476 51782 3528
rect 59722 3476 59728 3528
rect 59780 3516 59786 3528
rect 60737 3519 60795 3525
rect 60737 3516 60749 3519
rect 59780 3488 60749 3516
rect 59780 3476 59786 3488
rect 60737 3485 60749 3488
rect 60783 3485 60795 3519
rect 60737 3479 60795 3485
rect 61933 3519 61991 3525
rect 61933 3485 61945 3519
rect 61979 3485 61991 3519
rect 61933 3479 61991 3485
rect 25590 3408 25596 3460
rect 25648 3448 25654 3460
rect 43806 3448 43812 3460
rect 25648 3420 43812 3448
rect 25648 3408 25654 3420
rect 43806 3408 43812 3420
rect 43864 3408 43870 3460
rect 61948 3448 61976 3479
rect 65794 3476 65800 3528
rect 65852 3516 65858 3528
rect 66993 3519 67051 3525
rect 66993 3516 67005 3519
rect 65852 3488 67005 3516
rect 65852 3476 65858 3488
rect 66993 3485 67005 3488
rect 67039 3485 67051 3519
rect 66993 3479 67051 3485
rect 67358 3476 67364 3528
rect 67416 3516 67422 3528
rect 67453 3519 67511 3525
rect 67453 3516 67465 3519
rect 67416 3488 67465 3516
rect 67416 3476 67422 3488
rect 67453 3485 67465 3488
rect 67499 3485 67511 3519
rect 67453 3479 67511 3485
rect 62114 3448 62120 3460
rect 61948 3420 62120 3448
rect 62114 3408 62120 3420
rect 62172 3408 62178 3460
rect 22094 3380 22100 3392
rect 7668 3352 16574 3380
rect 22055 3352 22100 3380
rect 6825 3343 6883 3349
rect 22094 3340 22100 3352
rect 22152 3340 22158 3392
rect 24486 3340 24492 3392
rect 24544 3380 24550 3392
rect 26142 3380 26148 3392
rect 24544 3352 26148 3380
rect 24544 3340 24550 3352
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 44818 3340 44824 3392
rect 44876 3380 44882 3392
rect 45097 3383 45155 3389
rect 45097 3380 45109 3383
rect 44876 3352 45109 3380
rect 44876 3340 44882 3352
rect 45097 3349 45109 3352
rect 45143 3349 45155 3383
rect 60826 3380 60832 3392
rect 60787 3352 60832 3380
rect 45097 3343 45155 3349
rect 60826 3340 60832 3352
rect 60884 3340 60890 3392
rect 65978 3340 65984 3392
rect 66036 3380 66042 3392
rect 67545 3383 67603 3389
rect 67545 3380 67557 3383
rect 66036 3352 67557 3380
rect 66036 3340 66042 3352
rect 67545 3349 67557 3352
rect 67591 3349 67603 3383
rect 67545 3343 67603 3349
rect 1104 3290 68816 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 68816 3290
rect 1104 3216 68816 3238
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 37274 3176 37280 3188
rect 2004 3148 37280 3176
rect 2004 3136 2010 3148
rect 37274 3136 37280 3148
rect 37332 3136 37338 3188
rect 1762 3108 1768 3120
rect 1723 3080 1768 3108
rect 1762 3068 1768 3080
rect 1820 3068 1826 3120
rect 6822 3108 6828 3120
rect 6783 3080 6828 3108
rect 6822 3068 6828 3080
rect 6880 3068 6886 3120
rect 10594 3108 10600 3120
rect 10555 3080 10600 3108
rect 10594 3068 10600 3080
rect 10652 3068 10658 3120
rect 22094 3108 22100 3120
rect 22055 3080 22100 3108
rect 22094 3068 22100 3080
rect 22152 3068 22158 3120
rect 33505 3111 33563 3117
rect 33505 3077 33517 3111
rect 33551 3108 33563 3111
rect 34241 3111 34299 3117
rect 34241 3108 34253 3111
rect 33551 3080 34253 3108
rect 33551 3077 33563 3080
rect 33505 3071 33563 3077
rect 34241 3077 34253 3080
rect 34287 3077 34299 3111
rect 44818 3108 44824 3120
rect 44779 3080 44824 3108
rect 34241 3071 34299 3077
rect 44818 3068 44824 3080
rect 44876 3068 44882 3120
rect 60826 3108 60832 3120
rect 60787 3080 60832 3108
rect 60826 3068 60832 3080
rect 60884 3068 60890 3120
rect 65978 3108 65984 3120
rect 65939 3080 65984 3108
rect 65978 3068 65984 3080
rect 66036 3068 66042 3120
rect 1578 3040 1584 3052
rect 1539 3012 1584 3040
rect 1578 3000 1584 3012
rect 1636 3000 1642 3052
rect 3878 3040 3884 3052
rect 3839 3012 3884 3040
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 6638 3040 6644 3052
rect 6599 3012 6644 3040
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 10226 3040 10232 3052
rect 10139 3012 10232 3040
rect 10226 3000 10232 3012
rect 10284 3040 10290 3052
rect 10505 3043 10563 3049
rect 10505 3040 10517 3043
rect 10284 3012 10517 3040
rect 10284 3000 10290 3012
rect 10505 3009 10517 3012
rect 10551 3040 10563 3043
rect 19334 3040 19340 3052
rect 10551 3012 16574 3040
rect 19295 3012 19340 3040
rect 10551 3009 10563 3012
rect 10505 3003 10563 3009
rect 2774 2972 2780 2984
rect 2735 2944 2780 2972
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 3510 2932 3516 2984
rect 3568 2972 3574 2984
rect 4065 2975 4123 2981
rect 4065 2972 4077 2975
rect 3568 2944 4077 2972
rect 3568 2932 3574 2944
rect 4065 2941 4077 2944
rect 4111 2941 4123 2975
rect 4065 2935 4123 2941
rect 4341 2975 4399 2981
rect 4341 2941 4353 2975
rect 4387 2941 4399 2975
rect 7098 2972 7104 2984
rect 7059 2944 7104 2972
rect 4341 2935 4399 2941
rect 2866 2864 2872 2916
rect 2924 2904 2930 2916
rect 4356 2904 4384 2935
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 2924 2876 4384 2904
rect 2924 2864 2930 2876
rect 16546 2836 16574 3012
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 33410 3040 33416 3052
rect 33371 3012 33416 3040
rect 33410 3000 33416 3012
rect 33468 3000 33474 3052
rect 38102 3040 38108 3052
rect 38063 3012 38108 3040
rect 38102 3000 38108 3012
rect 38160 3000 38166 3052
rect 60642 3040 60648 3052
rect 60603 3012 60648 3040
rect 60642 3000 60648 3012
rect 60700 3000 60706 3052
rect 65794 3040 65800 3052
rect 65755 3012 65800 3040
rect 65794 3000 65800 3012
rect 65852 3000 65858 3052
rect 19518 2972 19524 2984
rect 19479 2944 19524 2972
rect 19518 2932 19524 2944
rect 19576 2932 19582 2984
rect 19978 2972 19984 2984
rect 19939 2944 19984 2972
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 21913 2975 21971 2981
rect 21913 2941 21925 2975
rect 21959 2972 21971 2975
rect 22738 2972 22744 2984
rect 21959 2944 22744 2972
rect 21959 2941 21971 2944
rect 21913 2935 21971 2941
rect 22738 2932 22744 2944
rect 22796 2932 22802 2984
rect 22833 2975 22891 2981
rect 22833 2941 22845 2975
rect 22879 2941 22891 2975
rect 22833 2935 22891 2941
rect 34057 2975 34115 2981
rect 34057 2941 34069 2975
rect 34103 2972 34115 2975
rect 34606 2972 34612 2984
rect 34103 2944 34612 2972
rect 34103 2941 34115 2944
rect 34057 2935 34115 2941
rect 22554 2864 22560 2916
rect 22612 2904 22618 2916
rect 22848 2904 22876 2935
rect 34606 2932 34612 2944
rect 34664 2932 34670 2984
rect 34790 2972 34796 2984
rect 34751 2944 34796 2972
rect 34790 2932 34796 2944
rect 34848 2932 34854 2984
rect 38286 2972 38292 2984
rect 38247 2944 38292 2972
rect 38286 2932 38292 2944
rect 38344 2932 38350 2984
rect 38654 2972 38660 2984
rect 38615 2944 38660 2972
rect 38654 2932 38660 2944
rect 38712 2932 38718 2984
rect 44177 2975 44235 2981
rect 44177 2941 44189 2975
rect 44223 2972 44235 2975
rect 44637 2975 44695 2981
rect 44637 2972 44649 2975
rect 44223 2944 44649 2972
rect 44223 2941 44235 2944
rect 44177 2935 44235 2941
rect 44637 2941 44649 2944
rect 44683 2941 44695 2975
rect 45094 2972 45100 2984
rect 45055 2944 45100 2972
rect 44637 2935 44695 2941
rect 45094 2932 45100 2944
rect 45152 2932 45158 2984
rect 61194 2972 61200 2984
rect 61155 2944 61200 2972
rect 61194 2932 61200 2944
rect 61252 2932 61258 2984
rect 67637 2975 67695 2981
rect 67637 2941 67649 2975
rect 67683 2972 67695 2975
rect 69566 2972 69572 2984
rect 67683 2944 69572 2972
rect 67683 2941 67695 2944
rect 67637 2935 67695 2941
rect 69566 2932 69572 2944
rect 69624 2932 69630 2984
rect 67082 2904 67088 2916
rect 22612 2876 22876 2904
rect 26206 2876 67088 2904
rect 22612 2864 22618 2876
rect 26206 2836 26234 2876
rect 67082 2864 67088 2876
rect 67140 2864 67146 2916
rect 16546 2808 26234 2836
rect 1104 2746 68816 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 68816 2746
rect 1104 2672 68816 2694
rect 2501 2635 2559 2641
rect 2501 2601 2513 2635
rect 2547 2632 2559 2635
rect 3510 2632 3516 2644
rect 2547 2604 3516 2632
rect 2547 2601 2559 2604
rect 2501 2595 2559 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 3970 2632 3976 2644
rect 3931 2604 3976 2632
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 10410 2592 10416 2644
rect 10468 2632 10474 2644
rect 10689 2635 10747 2641
rect 10689 2632 10701 2635
rect 10468 2604 10701 2632
rect 10468 2592 10474 2604
rect 10689 2601 10701 2604
rect 10735 2601 10747 2635
rect 17678 2632 17684 2644
rect 17639 2604 17684 2632
rect 10689 2595 10747 2601
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 19518 2632 19524 2644
rect 19479 2604 19524 2632
rect 19518 2592 19524 2604
rect 19576 2592 19582 2644
rect 22738 2632 22744 2644
rect 22699 2604 22744 2632
rect 22738 2592 22744 2604
rect 22796 2592 22802 2644
rect 32306 2632 32312 2644
rect 32267 2604 32312 2632
rect 32306 2592 32312 2604
rect 32364 2592 32370 2644
rect 34606 2592 34612 2644
rect 34664 2632 34670 2644
rect 34885 2635 34943 2641
rect 34885 2632 34897 2635
rect 34664 2604 34897 2632
rect 34664 2592 34670 2604
rect 34885 2601 34897 2604
rect 34931 2601 34943 2635
rect 34885 2595 34943 2601
rect 38197 2635 38255 2641
rect 38197 2601 38209 2635
rect 38243 2632 38255 2635
rect 38286 2632 38292 2644
rect 38243 2604 38292 2632
rect 38243 2601 38255 2604
rect 38197 2595 38255 2601
rect 38286 2592 38292 2604
rect 38344 2592 38350 2644
rect 46198 2592 46204 2644
rect 46256 2632 46262 2644
rect 46385 2635 46443 2641
rect 46385 2632 46397 2635
rect 46256 2604 46397 2632
rect 46256 2592 46262 2604
rect 46385 2601 46397 2604
rect 46431 2601 46443 2635
rect 62114 2632 62120 2644
rect 62075 2604 62120 2632
rect 46385 2595 46443 2601
rect 62114 2592 62120 2604
rect 62172 2592 62178 2644
rect 5810 2524 5816 2576
rect 5868 2564 5874 2576
rect 22005 2567 22063 2573
rect 5868 2536 6960 2564
rect 5868 2524 5874 2536
rect 6546 2496 6552 2508
rect 6507 2468 6552 2496
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 6932 2505 6960 2536
rect 22005 2533 22017 2567
rect 22051 2564 22063 2567
rect 25406 2564 25412 2576
rect 22051 2536 25412 2564
rect 22051 2533 22063 2536
rect 22005 2527 22063 2533
rect 25406 2524 25412 2536
rect 25464 2524 25470 2576
rect 25958 2524 25964 2576
rect 26016 2564 26022 2576
rect 43073 2567 43131 2573
rect 43073 2564 43085 2567
rect 26016 2536 43085 2564
rect 26016 2524 26022 2536
rect 43073 2533 43085 2536
rect 43119 2533 43131 2567
rect 43073 2527 43131 2533
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2465 6975 2499
rect 25314 2496 25320 2508
rect 6917 2459 6975 2465
rect 16546 2468 25320 2496
rect 2406 2428 2412 2440
rect 2367 2400 2412 2428
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3292 2400 3801 2428
rect 3292 2388 3298 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2428 5779 2431
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5767 2400 6377 2428
rect 5767 2397 5779 2400
rect 5721 2391 5779 2397
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 2424 2360 2452 2388
rect 16546 2360 16574 2468
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 19444 2437 19472 2468
rect 25314 2456 25320 2468
rect 25372 2496 25378 2508
rect 27430 2496 27436 2508
rect 25372 2468 27292 2496
rect 27391 2468 27436 2496
rect 25372 2456 25378 2468
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17460 2400 17509 2428
rect 17460 2388 17466 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 21324 2400 21833 2428
rect 21324 2388 21330 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27120 2400 27169 2428
rect 27120 2388 27126 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27264 2428 27292 2468
rect 27430 2456 27436 2468
rect 27488 2456 27494 2508
rect 33410 2496 33416 2508
rect 27540 2468 33416 2496
rect 27540 2428 27568 2468
rect 33410 2456 33416 2468
rect 33468 2456 33474 2508
rect 40604 2468 55214 2496
rect 27264 2400 27568 2428
rect 27157 2391 27215 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28445 2431 28503 2437
rect 28445 2428 28457 2431
rect 28408 2400 28457 2428
rect 28408 2388 28414 2400
rect 28445 2397 28457 2400
rect 28491 2397 28503 2431
rect 28445 2391 28503 2397
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 32493 2431 32551 2437
rect 32493 2428 32505 2431
rect 32272 2400 32505 2428
rect 32272 2388 32278 2400
rect 32493 2397 32505 2400
rect 32539 2397 32551 2431
rect 32493 2391 32551 2397
rect 37274 2388 37280 2440
rect 37332 2428 37338 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 37332 2400 38117 2428
rect 37332 2388 37338 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 2424 2332 16574 2360
rect 20898 2320 20904 2372
rect 20956 2360 20962 2372
rect 40604 2360 40632 2468
rect 20956 2332 40632 2360
rect 40696 2400 43024 2428
rect 20956 2320 20962 2332
rect 20806 2252 20812 2304
rect 20864 2292 20870 2304
rect 28629 2295 28687 2301
rect 28629 2292 28641 2295
rect 20864 2264 28641 2292
rect 20864 2252 20870 2264
rect 28629 2261 28641 2264
rect 28675 2261 28687 2295
rect 28629 2255 28687 2261
rect 32122 2252 32128 2304
rect 32180 2292 32186 2304
rect 40696 2292 40724 2400
rect 42518 2320 42524 2372
rect 42576 2360 42582 2372
rect 42889 2363 42947 2369
rect 42889 2360 42901 2363
rect 42576 2332 42901 2360
rect 42576 2320 42582 2332
rect 42889 2329 42901 2332
rect 42935 2329 42947 2363
rect 42996 2360 43024 2400
rect 55186 2360 55214 2468
rect 56042 2388 56048 2440
rect 56100 2428 56106 2440
rect 56137 2431 56195 2437
rect 56137 2428 56149 2431
rect 56100 2400 56149 2428
rect 56100 2388 56106 2400
rect 56137 2397 56149 2400
rect 56183 2397 56195 2431
rect 56137 2391 56195 2397
rect 56336 2400 58020 2428
rect 56336 2360 56364 2400
rect 42996 2332 45554 2360
rect 55186 2332 56364 2360
rect 42889 2323 42947 2329
rect 32180 2264 40724 2292
rect 45526 2292 45554 2332
rect 56410 2320 56416 2372
rect 56468 2360 56474 2372
rect 57992 2360 58020 2400
rect 65058 2388 65064 2440
rect 65116 2428 65122 2440
rect 65613 2431 65671 2437
rect 65613 2428 65625 2431
rect 65116 2400 65625 2428
rect 65116 2388 65122 2400
rect 65613 2397 65625 2400
rect 65659 2397 65671 2431
rect 65613 2391 65671 2397
rect 65889 2363 65947 2369
rect 65889 2360 65901 2363
rect 56468 2332 56513 2360
rect 57992 2332 65901 2360
rect 56468 2320 56474 2332
rect 65889 2329 65901 2332
rect 65935 2329 65947 2363
rect 65889 2323 65947 2329
rect 67269 2363 67327 2369
rect 67269 2329 67281 2363
rect 67315 2360 67327 2363
rect 67634 2360 67640 2372
rect 67315 2332 67640 2360
rect 67315 2329 67327 2332
rect 67269 2323 67327 2329
rect 67634 2320 67640 2332
rect 67692 2320 67698 2372
rect 67361 2295 67419 2301
rect 67361 2292 67373 2295
rect 45526 2264 67373 2292
rect 32180 2252 32186 2264
rect 67361 2261 67373 2264
rect 67407 2261 67419 2295
rect 67361 2255 67419 2261
rect 1104 2202 68816 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 68816 2202
rect 1104 2128 68816 2150
rect 26602 1980 26608 2032
rect 26660 2020 26666 2032
rect 56410 2020 56416 2032
rect 26660 1992 56416 2020
rect 26660 1980 26666 1992
rect 56410 1980 56416 1992
rect 56468 1980 56474 2032
rect 50614 1300 50620 1352
rect 50672 1340 50678 1352
rect 66162 1340 66168 1352
rect 50672 1312 66168 1340
rect 50672 1300 50678 1312
rect 66162 1300 66168 1312
rect 66220 1300 66226 1352
<< via1 >>
rect 19574 69606 19626 69658
rect 19638 69606 19690 69658
rect 19702 69606 19754 69658
rect 19766 69606 19818 69658
rect 19830 69606 19882 69658
rect 50294 69606 50346 69658
rect 50358 69606 50410 69658
rect 50422 69606 50474 69658
rect 50486 69606 50538 69658
rect 50550 69606 50602 69658
rect 14188 69436 14240 69488
rect 19340 69436 19392 69488
rect 20628 69436 20680 69488
rect 35624 69479 35676 69488
rect 35624 69445 35633 69479
rect 35633 69445 35667 69479
rect 35667 69445 35676 69479
rect 35624 69436 35676 69445
rect 68284 69436 68336 69488
rect 1400 69411 1452 69420
rect 1400 69377 1409 69411
rect 1409 69377 1443 69411
rect 1443 69377 1452 69411
rect 1400 69368 1452 69377
rect 7748 69368 7800 69420
rect 46480 69368 46532 69420
rect 1584 69343 1636 69352
rect 1584 69309 1593 69343
rect 1593 69309 1627 69343
rect 1627 69309 1636 69343
rect 1584 69300 1636 69309
rect 55404 69368 55456 69420
rect 57244 69368 57296 69420
rect 59728 69300 59780 69352
rect 65064 69300 65116 69352
rect 66352 69300 66404 69352
rect 14832 69232 14884 69284
rect 20260 69232 20312 69284
rect 21640 69232 21692 69284
rect 36912 69232 36964 69284
rect 2504 69207 2556 69216
rect 2504 69173 2513 69207
rect 2513 69173 2547 69207
rect 2547 69173 2556 69207
rect 2504 69164 2556 69173
rect 4804 69207 4856 69216
rect 4804 69173 4813 69207
rect 4813 69173 4847 69207
rect 4847 69173 4856 69207
rect 4804 69164 4856 69173
rect 6000 69164 6052 69216
rect 8024 69207 8076 69216
rect 8024 69173 8033 69207
rect 8033 69173 8067 69207
rect 8067 69173 8076 69207
rect 8024 69164 8076 69173
rect 11704 69207 11756 69216
rect 11704 69173 11713 69207
rect 11713 69173 11747 69207
rect 11747 69173 11756 69207
rect 11704 69164 11756 69173
rect 16856 69207 16908 69216
rect 16856 69173 16865 69207
rect 16865 69173 16899 69207
rect 16899 69173 16908 69207
rect 16856 69164 16908 69173
rect 24860 69207 24912 69216
rect 24860 69173 24869 69207
rect 24869 69173 24903 69207
rect 24903 69173 24912 69207
rect 24860 69164 24912 69173
rect 27344 69207 27396 69216
rect 27344 69173 27353 69207
rect 27353 69173 27387 69207
rect 27387 69173 27396 69207
rect 27344 69164 27396 69173
rect 31208 69207 31260 69216
rect 31208 69173 31217 69207
rect 31217 69173 31251 69207
rect 31251 69173 31260 69207
rect 31208 69164 31260 69173
rect 36636 69207 36688 69216
rect 36636 69173 36645 69207
rect 36645 69173 36679 69207
rect 36679 69173 36688 69207
rect 36636 69164 36688 69173
rect 37280 69164 37332 69216
rect 39028 69207 39080 69216
rect 39028 69173 39037 69207
rect 39037 69173 39071 69207
rect 39071 69173 39080 69207
rect 39028 69164 39080 69173
rect 41420 69207 41472 69216
rect 41420 69173 41429 69207
rect 41429 69173 41463 69207
rect 41463 69173 41472 69207
rect 41420 69164 41472 69173
rect 42892 69207 42944 69216
rect 42892 69173 42901 69207
rect 42901 69173 42935 69207
rect 42935 69173 42944 69207
rect 42892 69164 42944 69173
rect 45192 69164 45244 69216
rect 46112 69207 46164 69216
rect 46112 69173 46121 69207
rect 46121 69173 46155 69207
rect 46155 69173 46164 69207
rect 46112 69164 46164 69173
rect 46572 69164 46624 69216
rect 50712 69207 50764 69216
rect 50712 69173 50721 69207
rect 50721 69173 50755 69207
rect 50755 69173 50764 69207
rect 50712 69164 50764 69173
rect 52920 69207 52972 69216
rect 52920 69173 52929 69207
rect 52929 69173 52963 69207
rect 52963 69173 52972 69207
rect 52920 69164 52972 69173
rect 55680 69207 55732 69216
rect 55680 69173 55689 69207
rect 55689 69173 55723 69207
rect 55723 69173 55732 69207
rect 55680 69164 55732 69173
rect 56508 69207 56560 69216
rect 56508 69173 56517 69207
rect 56517 69173 56551 69207
rect 56551 69173 56560 69207
rect 56508 69164 56560 69173
rect 57336 69207 57388 69216
rect 57336 69173 57345 69207
rect 57345 69173 57379 69207
rect 57379 69173 57388 69207
rect 57336 69164 57388 69173
rect 58072 69164 58124 69216
rect 60648 69207 60700 69216
rect 60648 69173 60657 69207
rect 60657 69173 60691 69207
rect 60691 69173 60700 69207
rect 60648 69164 60700 69173
rect 62212 69207 62264 69216
rect 62212 69173 62221 69207
rect 62221 69173 62255 69207
rect 62255 69173 62264 69207
rect 62212 69164 62264 69173
rect 64972 69164 65024 69216
rect 66260 69164 66312 69216
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 34934 69062 34986 69114
rect 34998 69062 35050 69114
rect 35062 69062 35114 69114
rect 35126 69062 35178 69114
rect 35190 69062 35242 69114
rect 65654 69062 65706 69114
rect 65718 69062 65770 69114
rect 65782 69062 65834 69114
rect 65846 69062 65898 69114
rect 65910 69062 65962 69114
rect 11612 68892 11664 68944
rect 2504 68824 2556 68876
rect 2780 68867 2832 68876
rect 2780 68833 2789 68867
rect 2789 68833 2823 68867
rect 2823 68833 2832 68867
rect 2780 68824 2832 68833
rect 6000 68867 6052 68876
rect 6000 68833 6009 68867
rect 6009 68833 6043 68867
rect 6043 68833 6052 68867
rect 6000 68824 6052 68833
rect 6460 68867 6512 68876
rect 6460 68833 6469 68867
rect 6469 68833 6503 68867
rect 6503 68833 6512 68867
rect 6460 68824 6512 68833
rect 11704 68824 11756 68876
rect 16764 68892 16816 68944
rect 16856 68824 16908 68876
rect 52828 68892 52880 68944
rect 24860 68824 24912 68876
rect 25136 68867 25188 68876
rect 25136 68833 25145 68867
rect 25145 68833 25179 68867
rect 25179 68833 25188 68867
rect 25136 68824 25188 68833
rect 27344 68824 27396 68876
rect 27712 68867 27764 68876
rect 27712 68833 27721 68867
rect 27721 68833 27755 68867
rect 27755 68833 27764 68867
rect 27712 68824 27764 68833
rect 31208 68824 31260 68876
rect 31576 68824 31628 68876
rect 36636 68824 36688 68876
rect 36728 68867 36780 68876
rect 36728 68833 36737 68867
rect 36737 68833 36771 68867
rect 36771 68833 36780 68867
rect 36728 68824 36780 68833
rect 41420 68824 41472 68876
rect 41880 68867 41932 68876
rect 41880 68833 41889 68867
rect 41889 68833 41923 68867
rect 41923 68833 41932 68867
rect 41880 68824 41932 68833
rect 42892 68824 42944 68876
rect 43168 68867 43220 68876
rect 43168 68833 43177 68867
rect 43177 68833 43211 68867
rect 43211 68833 43220 68867
rect 43168 68824 43220 68833
rect 46112 68824 46164 68876
rect 46572 68867 46624 68876
rect 46572 68833 46581 68867
rect 46581 68833 46615 68867
rect 46615 68833 46624 68867
rect 46572 68824 46624 68833
rect 47032 68867 47084 68876
rect 47032 68833 47041 68867
rect 47041 68833 47075 68867
rect 47075 68833 47084 68867
rect 47032 68824 47084 68833
rect 50712 68824 50764 68876
rect 51540 68867 51592 68876
rect 51540 68833 51549 68867
rect 51549 68833 51583 68867
rect 51583 68833 51592 68867
rect 51540 68824 51592 68833
rect 52920 68824 52972 68876
rect 60556 68892 60608 68944
rect 56508 68824 56560 68876
rect 56692 68867 56744 68876
rect 56692 68833 56701 68867
rect 56701 68833 56735 68867
rect 56735 68833 56744 68867
rect 56692 68824 56744 68833
rect 60648 68824 60700 68876
rect 62212 68824 62264 68876
rect 63132 68824 63184 68876
rect 66260 68867 66312 68876
rect 66260 68833 66269 68867
rect 66269 68833 66303 68867
rect 66303 68833 66312 68867
rect 66260 68824 66312 68833
rect 69572 68824 69624 68876
rect 4620 68799 4672 68808
rect 4620 68765 4629 68799
rect 4629 68765 4663 68799
rect 4663 68765 4672 68799
rect 4620 68756 4672 68765
rect 5908 68756 5960 68808
rect 10416 68799 10468 68808
rect 10416 68765 10425 68799
rect 10425 68765 10459 68799
rect 10459 68765 10468 68799
rect 10416 68756 10468 68765
rect 15476 68799 15528 68808
rect 15476 68765 15485 68799
rect 15485 68765 15519 68799
rect 15519 68765 15528 68799
rect 15476 68756 15528 68765
rect 38936 68799 38988 68808
rect 38936 68765 38945 68799
rect 38945 68765 38979 68799
rect 38979 68765 38988 68799
rect 38936 68756 38988 68765
rect 39856 68756 39908 68808
rect 1860 68688 1912 68740
rect 24860 68731 24912 68740
rect 24860 68697 24869 68731
rect 24869 68697 24903 68731
rect 24903 68697 24912 68731
rect 24860 68688 24912 68697
rect 27252 68731 27304 68740
rect 27252 68697 27261 68731
rect 27261 68697 27295 68731
rect 27295 68697 27304 68731
rect 27252 68688 27304 68697
rect 31208 68731 31260 68740
rect 31208 68697 31217 68731
rect 31217 68697 31251 68731
rect 31251 68697 31260 68731
rect 31208 68688 31260 68697
rect 36544 68688 36596 68740
rect 41420 68688 41472 68740
rect 42800 68731 42852 68740
rect 42800 68697 42809 68731
rect 42809 68697 42843 68731
rect 42843 68697 42852 68731
rect 42800 68688 42852 68697
rect 4712 68663 4764 68672
rect 4712 68629 4721 68663
rect 4721 68629 4755 68663
rect 4755 68629 4764 68663
rect 4712 68620 4764 68629
rect 15476 68620 15528 68672
rect 27160 68620 27212 68672
rect 39764 68620 39816 68672
rect 42616 68620 42668 68672
rect 48964 68799 49016 68808
rect 48964 68765 48973 68799
rect 48973 68765 49007 68799
rect 49007 68765 49016 68799
rect 48964 68756 49016 68765
rect 59728 68799 59780 68808
rect 59728 68765 59737 68799
rect 59737 68765 59771 68799
rect 59771 68765 59780 68799
rect 59728 68756 59780 68765
rect 52920 68731 52972 68740
rect 52920 68697 52929 68731
rect 52929 68697 52963 68731
rect 52963 68697 52972 68731
rect 52920 68688 52972 68697
rect 56416 68731 56468 68740
rect 56416 68697 56425 68731
rect 56425 68697 56459 68731
rect 56459 68697 56468 68731
rect 56416 68688 56468 68697
rect 62948 68731 63000 68740
rect 62948 68697 62957 68731
rect 62957 68697 62991 68731
rect 62991 68697 63000 68731
rect 62948 68688 63000 68697
rect 45376 68663 45428 68672
rect 45376 68629 45385 68663
rect 45385 68629 45419 68663
rect 45419 68629 45428 68663
rect 45376 68620 45428 68629
rect 59728 68620 59780 68672
rect 67088 68688 67140 68740
rect 65708 68663 65760 68672
rect 65708 68629 65717 68663
rect 65717 68629 65751 68663
rect 65751 68629 65760 68663
rect 65708 68620 65760 68629
rect 19574 68518 19626 68570
rect 19638 68518 19690 68570
rect 19702 68518 19754 68570
rect 19766 68518 19818 68570
rect 19830 68518 19882 68570
rect 50294 68518 50346 68570
rect 50358 68518 50410 68570
rect 50422 68518 50474 68570
rect 50486 68518 50538 68570
rect 50550 68518 50602 68570
rect 1860 68459 1912 68468
rect 1860 68425 1869 68459
rect 1869 68425 1903 68459
rect 1903 68425 1912 68459
rect 1860 68416 1912 68425
rect 4620 68416 4672 68468
rect 23296 68416 23348 68468
rect 24860 68416 24912 68468
rect 27252 68459 27304 68468
rect 27252 68425 27261 68459
rect 27261 68425 27295 68459
rect 27295 68425 27304 68459
rect 27252 68416 27304 68425
rect 31208 68416 31260 68468
rect 36544 68459 36596 68468
rect 36544 68425 36553 68459
rect 36553 68425 36587 68459
rect 36587 68425 36596 68459
rect 36544 68416 36596 68425
rect 42616 68416 42668 68468
rect 42800 68459 42852 68468
rect 42800 68425 42809 68459
rect 42809 68425 42843 68459
rect 42843 68425 42852 68459
rect 42800 68416 42852 68425
rect 39764 68391 39816 68400
rect 2044 68280 2096 68332
rect 24676 68323 24728 68332
rect 24676 68289 24685 68323
rect 24685 68289 24719 68323
rect 24719 68289 24728 68323
rect 24676 68280 24728 68289
rect 27160 68323 27212 68332
rect 27160 68289 27169 68323
rect 27169 68289 27203 68323
rect 27203 68289 27212 68323
rect 39764 68357 39773 68391
rect 39773 68357 39807 68391
rect 39807 68357 39816 68391
rect 39764 68348 39816 68357
rect 39856 68348 39908 68400
rect 45376 68391 45428 68400
rect 45376 68357 45385 68391
rect 45385 68357 45419 68391
rect 45419 68357 45428 68391
rect 45376 68348 45428 68357
rect 52920 68416 52972 68468
rect 56416 68416 56468 68468
rect 62948 68416 63000 68468
rect 57244 68348 57296 68400
rect 58072 68391 58124 68400
rect 58072 68357 58081 68391
rect 58081 68357 58115 68391
rect 58115 68357 58124 68391
rect 58072 68348 58124 68357
rect 65708 68391 65760 68400
rect 65708 68357 65717 68391
rect 65717 68357 65751 68391
rect 65751 68357 65760 68391
rect 65708 68348 65760 68357
rect 31024 68323 31076 68332
rect 27160 68280 27212 68289
rect 31024 68289 31033 68323
rect 31033 68289 31067 68323
rect 31067 68289 31076 68323
rect 31024 68280 31076 68289
rect 36452 68323 36504 68332
rect 36452 68289 36461 68323
rect 36461 68289 36495 68323
rect 36495 68289 36504 68323
rect 36452 68280 36504 68289
rect 37280 68323 37332 68332
rect 37280 68289 37289 68323
rect 37289 68289 37323 68323
rect 37323 68289 37332 68323
rect 37280 68280 37332 68289
rect 39028 68280 39080 68332
rect 45192 68323 45244 68332
rect 3056 68212 3108 68264
rect 3332 68255 3384 68264
rect 3332 68221 3341 68255
rect 3341 68221 3375 68255
rect 3375 68221 3384 68255
rect 3332 68212 3384 68221
rect 37556 68212 37608 68264
rect 38016 68255 38068 68264
rect 38016 68221 38025 68255
rect 38025 68221 38059 68255
rect 38059 68221 38068 68255
rect 38016 68212 38068 68221
rect 39304 68212 39356 68264
rect 45192 68289 45201 68323
rect 45201 68289 45235 68323
rect 45235 68289 45244 68323
rect 45192 68280 45244 68289
rect 48964 68280 49016 68332
rect 52736 68323 52788 68332
rect 52736 68289 52745 68323
rect 52745 68289 52779 68323
rect 52779 68289 52788 68323
rect 52736 68280 52788 68289
rect 56232 68323 56284 68332
rect 56232 68289 56241 68323
rect 56241 68289 56275 68323
rect 56275 68289 56284 68323
rect 56232 68280 56284 68289
rect 45744 68255 45796 68264
rect 45744 68221 45753 68255
rect 45753 68221 45787 68255
rect 45787 68221 45796 68255
rect 45744 68212 45796 68221
rect 50252 68212 50304 68264
rect 42708 68144 42760 68196
rect 50160 68144 50212 68196
rect 57336 68280 57388 68332
rect 61568 68323 61620 68332
rect 61568 68289 61577 68323
rect 61577 68289 61611 68323
rect 61611 68289 61620 68323
rect 61568 68280 61620 68289
rect 64972 68280 65024 68332
rect 58072 68212 58124 68264
rect 65064 68255 65116 68264
rect 65064 68221 65073 68255
rect 65073 68221 65107 68255
rect 65107 68221 65116 68255
rect 65064 68212 65116 68221
rect 66996 68255 67048 68264
rect 66996 68221 67005 68255
rect 67005 68221 67039 68255
rect 67039 68221 67048 68255
rect 66996 68212 67048 68221
rect 67272 68144 67324 68196
rect 29184 68076 29236 68128
rect 30288 68076 30340 68128
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 34934 67974 34986 68026
rect 34998 67974 35050 68026
rect 35062 67974 35114 68026
rect 35126 67974 35178 68026
rect 35190 67974 35242 68026
rect 65654 67974 65706 68026
rect 65718 67974 65770 68026
rect 65782 67974 65834 68026
rect 65846 67974 65898 68026
rect 65910 67974 65962 68026
rect 37556 67915 37608 67924
rect 37556 67881 37565 67915
rect 37565 67881 37599 67915
rect 37599 67881 37608 67915
rect 37556 67872 37608 67881
rect 41420 67915 41472 67924
rect 41420 67881 41429 67915
rect 41429 67881 41463 67915
rect 41463 67881 41472 67915
rect 41420 67872 41472 67881
rect 50252 67915 50304 67924
rect 50252 67881 50261 67915
rect 50261 67881 50295 67915
rect 50295 67881 50304 67915
rect 50252 67872 50304 67881
rect 66352 67872 66404 67924
rect 67088 67915 67140 67924
rect 67088 67881 67097 67915
rect 67097 67881 67131 67915
rect 67131 67881 67140 67915
rect 67088 67872 67140 67881
rect 2320 67779 2372 67788
rect 2320 67745 2329 67779
rect 2329 67745 2363 67779
rect 2363 67745 2372 67779
rect 2320 67736 2372 67745
rect 4804 67804 4856 67856
rect 4712 67779 4764 67788
rect 4712 67745 4721 67779
rect 4721 67745 4755 67779
rect 4755 67745 4764 67779
rect 4712 67736 4764 67745
rect 5172 67779 5224 67788
rect 5172 67745 5181 67779
rect 5181 67745 5215 67779
rect 5215 67745 5224 67779
rect 5172 67736 5224 67745
rect 2044 67711 2096 67720
rect 2044 67677 2053 67711
rect 2053 67677 2087 67711
rect 2087 67677 2096 67711
rect 2044 67668 2096 67677
rect 2320 67600 2372 67652
rect 24676 67736 24728 67788
rect 31024 67736 31076 67788
rect 37464 67711 37516 67720
rect 37464 67677 37473 67711
rect 37473 67677 37507 67711
rect 37507 67677 37516 67711
rect 37464 67668 37516 67677
rect 41328 67711 41380 67720
rect 41328 67677 41337 67711
rect 41337 67677 41371 67711
rect 41371 67677 41380 67711
rect 41328 67668 41380 67677
rect 50160 67711 50212 67720
rect 50160 67677 50169 67711
rect 50169 67677 50203 67711
rect 50203 67677 50212 67711
rect 50160 67668 50212 67677
rect 66720 67668 66772 67720
rect 67732 67711 67784 67720
rect 67732 67677 67741 67711
rect 67741 67677 67775 67711
rect 67775 67677 67784 67711
rect 67732 67668 67784 67677
rect 38568 67600 38620 67652
rect 19574 67430 19626 67482
rect 19638 67430 19690 67482
rect 19702 67430 19754 67482
rect 19766 67430 19818 67482
rect 19830 67430 19882 67482
rect 50294 67430 50346 67482
rect 50358 67430 50410 67482
rect 50422 67430 50474 67482
rect 50486 67430 50538 67482
rect 50550 67430 50602 67482
rect 67640 67303 67692 67312
rect 67640 67269 67649 67303
rect 67649 67269 67683 67303
rect 67683 67269 67692 67303
rect 67640 67260 67692 67269
rect 1584 67235 1636 67244
rect 1584 67201 1593 67235
rect 1593 67201 1627 67235
rect 1627 67201 1636 67235
rect 1584 67192 1636 67201
rect 2044 67192 2096 67244
rect 2596 67192 2648 67244
rect 2872 67124 2924 67176
rect 3056 67167 3108 67176
rect 3056 67133 3065 67167
rect 3065 67133 3099 67167
rect 3099 67133 3108 67167
rect 3056 67124 3108 67133
rect 5172 67167 5224 67176
rect 5172 67133 5181 67167
rect 5181 67133 5215 67167
rect 5215 67133 5224 67167
rect 5172 67124 5224 67133
rect 40960 67124 41012 67176
rect 41328 67124 41380 67176
rect 36452 67056 36504 67108
rect 37004 67056 37056 67108
rect 67548 67124 67600 67176
rect 66996 67056 67048 67108
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 34934 66886 34986 66938
rect 34998 66886 35050 66938
rect 35062 66886 35114 66938
rect 35126 66886 35178 66938
rect 35190 66886 35242 66938
rect 65654 66886 65706 66938
rect 65718 66886 65770 66938
rect 65782 66886 65834 66938
rect 65846 66886 65898 66938
rect 65910 66886 65962 66938
rect 66996 66827 67048 66836
rect 66996 66793 67005 66827
rect 67005 66793 67039 66827
rect 67039 66793 67048 66827
rect 66996 66784 67048 66793
rect 67548 66827 67600 66836
rect 67548 66793 67557 66827
rect 67557 66793 67591 66827
rect 67591 66793 67600 66827
rect 67548 66784 67600 66793
rect 2780 66691 2832 66700
rect 2780 66657 2789 66691
rect 2789 66657 2823 66691
rect 2823 66657 2832 66691
rect 2780 66648 2832 66657
rect 5908 66648 5960 66700
rect 10416 66648 10468 66700
rect 1400 66623 1452 66632
rect 1400 66589 1409 66623
rect 1409 66589 1443 66623
rect 1443 66589 1452 66623
rect 1400 66580 1452 66589
rect 4068 66580 4120 66632
rect 50160 66580 50212 66632
rect 67456 66623 67508 66632
rect 67456 66589 67465 66623
rect 67465 66589 67499 66623
rect 67499 66589 67508 66623
rect 67456 66580 67508 66589
rect 1584 66555 1636 66564
rect 1584 66521 1593 66555
rect 1593 66521 1627 66555
rect 1627 66521 1636 66555
rect 1584 66512 1636 66521
rect 4712 66444 4764 66496
rect 37464 66444 37516 66496
rect 19574 66342 19626 66394
rect 19638 66342 19690 66394
rect 19702 66342 19754 66394
rect 19766 66342 19818 66394
rect 19830 66342 19882 66394
rect 50294 66342 50346 66394
rect 50358 66342 50410 66394
rect 50422 66342 50474 66394
rect 50486 66342 50538 66394
rect 50550 66342 50602 66394
rect 1584 66240 1636 66292
rect 2596 66147 2648 66156
rect 2596 66113 2605 66147
rect 2605 66113 2639 66147
rect 2639 66113 2648 66147
rect 2596 66104 2648 66113
rect 4068 66104 4120 66156
rect 25136 66104 25188 66156
rect 36084 66147 36136 66156
rect 36084 66113 36093 66147
rect 36093 66113 36127 66147
rect 36127 66113 36136 66147
rect 36084 66104 36136 66113
rect 3424 65968 3476 66020
rect 5264 66036 5316 66088
rect 52736 66104 52788 66156
rect 53104 66104 53156 66156
rect 36360 66079 36412 66088
rect 36360 66045 36369 66079
rect 36369 66045 36403 66079
rect 36403 66045 36412 66079
rect 36360 66036 36412 66045
rect 46480 65968 46532 66020
rect 67364 66036 67416 66088
rect 67548 66079 67600 66088
rect 67548 66045 67557 66079
rect 67557 66045 67591 66079
rect 67591 66045 67600 66079
rect 67548 66036 67600 66045
rect 66996 65968 67048 66020
rect 35900 65943 35952 65952
rect 35900 65909 35909 65943
rect 35909 65909 35943 65943
rect 35943 65909 35952 65943
rect 35900 65900 35952 65909
rect 36360 65900 36412 65952
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 34934 65798 34986 65850
rect 34998 65798 35050 65850
rect 35062 65798 35114 65850
rect 35126 65798 35178 65850
rect 35190 65798 35242 65850
rect 65654 65798 65706 65850
rect 65718 65798 65770 65850
rect 65782 65798 65834 65850
rect 65846 65798 65898 65850
rect 65910 65798 65962 65850
rect 66996 65739 67048 65748
rect 66996 65705 67005 65739
rect 67005 65705 67039 65739
rect 67039 65705 67048 65739
rect 66996 65696 67048 65705
rect 67364 65696 67416 65748
rect 1768 65492 1820 65544
rect 2872 65467 2924 65476
rect 2872 65433 2881 65467
rect 2881 65433 2915 65467
rect 2915 65433 2924 65467
rect 2872 65424 2924 65433
rect 4068 65492 4120 65544
rect 33968 65492 34020 65544
rect 35900 65492 35952 65544
rect 67272 65492 67324 65544
rect 4344 65424 4396 65476
rect 4804 65467 4856 65476
rect 4804 65433 4813 65467
rect 4813 65433 4847 65467
rect 4847 65433 4856 65467
rect 4804 65424 4856 65433
rect 1952 65356 2004 65408
rect 23112 65356 23164 65408
rect 36268 65356 36320 65408
rect 19574 65254 19626 65306
rect 19638 65254 19690 65306
rect 19702 65254 19754 65306
rect 19766 65254 19818 65306
rect 19830 65254 19882 65306
rect 50294 65254 50346 65306
rect 50358 65254 50410 65306
rect 50422 65254 50474 65306
rect 50486 65254 50538 65306
rect 50550 65254 50602 65306
rect 4804 65152 4856 65204
rect 50160 65152 50212 65204
rect 1952 65127 2004 65136
rect 1952 65093 1961 65127
rect 1961 65093 1995 65127
rect 1995 65093 2004 65127
rect 1952 65084 2004 65093
rect 1768 65059 1820 65068
rect 1768 65025 1777 65059
rect 1777 65025 1811 65059
rect 1811 65025 1820 65059
rect 1768 65016 1820 65025
rect 4068 65059 4120 65068
rect 4068 65025 4077 65059
rect 4077 65025 4111 65059
rect 4111 65025 4120 65059
rect 4068 65016 4120 65025
rect 36084 65059 36136 65068
rect 36084 65025 36093 65059
rect 36093 65025 36127 65059
rect 36127 65025 36136 65059
rect 36084 65016 36136 65025
rect 36268 65059 36320 65068
rect 36268 65025 36277 65059
rect 36277 65025 36311 65059
rect 36311 65025 36320 65059
rect 36268 65016 36320 65025
rect 36360 65059 36412 65068
rect 36360 65025 36369 65059
rect 36369 65025 36403 65059
rect 36403 65025 36412 65059
rect 38292 65059 38344 65068
rect 36360 65016 36412 65025
rect 38292 65025 38301 65059
rect 38301 65025 38335 65059
rect 38335 65025 38344 65059
rect 38292 65016 38344 65025
rect 3608 64991 3660 65000
rect 3608 64957 3617 64991
rect 3617 64957 3651 64991
rect 3651 64957 3660 64991
rect 3608 64948 3660 64957
rect 4344 64991 4396 65000
rect 4344 64957 4353 64991
rect 4353 64957 4387 64991
rect 4387 64957 4396 64991
rect 4344 64948 4396 64957
rect 15476 64948 15528 65000
rect 36544 64948 36596 65000
rect 38200 64812 38252 64864
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 34934 64710 34986 64762
rect 34998 64710 35050 64762
rect 35062 64710 35114 64762
rect 35126 64710 35178 64762
rect 35190 64710 35242 64762
rect 65654 64710 65706 64762
rect 65718 64710 65770 64762
rect 65782 64710 65834 64762
rect 65846 64710 65898 64762
rect 65910 64710 65962 64762
rect 1400 64608 1452 64660
rect 36360 64540 36412 64592
rect 36728 64540 36780 64592
rect 36636 64404 36688 64456
rect 38292 64608 38344 64660
rect 38200 64447 38252 64456
rect 38200 64413 38234 64447
rect 38234 64413 38252 64447
rect 38200 64404 38252 64413
rect 36544 64336 36596 64388
rect 38108 64336 38160 64388
rect 37280 64311 37332 64320
rect 37280 64277 37289 64311
rect 37289 64277 37323 64311
rect 37323 64277 37332 64311
rect 37280 64268 37332 64277
rect 37740 64268 37792 64320
rect 19574 64166 19626 64218
rect 19638 64166 19690 64218
rect 19702 64166 19754 64218
rect 19766 64166 19818 64218
rect 19830 64166 19882 64218
rect 50294 64166 50346 64218
rect 50358 64166 50410 64218
rect 50422 64166 50474 64218
rect 50486 64166 50538 64218
rect 50550 64166 50602 64218
rect 36728 64107 36780 64116
rect 36728 64073 36737 64107
rect 36737 64073 36771 64107
rect 36771 64073 36780 64107
rect 36728 64064 36780 64073
rect 37280 64064 37332 64116
rect 38016 64064 38068 64116
rect 34704 63928 34756 63980
rect 37648 63996 37700 64048
rect 36820 63928 36872 63980
rect 37740 63971 37792 63980
rect 37740 63937 37749 63971
rect 37749 63937 37783 63971
rect 37783 63937 37792 63971
rect 37740 63928 37792 63937
rect 33416 63860 33468 63912
rect 33968 63903 34020 63912
rect 33968 63869 33977 63903
rect 33977 63869 34011 63903
rect 34011 63869 34020 63903
rect 33968 63860 34020 63869
rect 37648 63860 37700 63912
rect 35348 63767 35400 63776
rect 35348 63733 35357 63767
rect 35357 63733 35391 63767
rect 35391 63733 35400 63767
rect 35348 63724 35400 63733
rect 37280 63724 37332 63776
rect 66260 63724 66312 63776
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 34934 63622 34986 63674
rect 34998 63622 35050 63674
rect 35062 63622 35114 63674
rect 35126 63622 35178 63674
rect 35190 63622 35242 63674
rect 65654 63622 65706 63674
rect 65718 63622 65770 63674
rect 65782 63622 65834 63674
rect 65846 63622 65898 63674
rect 65910 63622 65962 63674
rect 34704 63563 34756 63572
rect 34704 63529 34713 63563
rect 34713 63529 34747 63563
rect 34747 63529 34756 63563
rect 34704 63520 34756 63529
rect 35808 63520 35860 63572
rect 36084 63520 36136 63572
rect 36636 63520 36688 63572
rect 25320 63452 25372 63504
rect 61568 63452 61620 63504
rect 35348 63384 35400 63436
rect 36452 63384 36504 63436
rect 37280 63384 37332 63436
rect 38016 63384 38068 63436
rect 66260 63427 66312 63436
rect 66260 63393 66269 63427
rect 66269 63393 66303 63427
rect 66303 63393 66312 63427
rect 66260 63384 66312 63393
rect 1400 63359 1452 63368
rect 1400 63325 1409 63359
rect 1409 63325 1443 63359
rect 1443 63325 1452 63359
rect 1400 63316 1452 63325
rect 24400 63316 24452 63368
rect 24860 63291 24912 63300
rect 24860 63257 24869 63291
rect 24869 63257 24903 63291
rect 24903 63257 24912 63291
rect 24860 63248 24912 63257
rect 35716 63316 35768 63368
rect 36820 63316 36872 63368
rect 31944 63180 31996 63232
rect 36084 63180 36136 63232
rect 36636 63248 36688 63300
rect 37740 63316 37792 63368
rect 68100 63359 68152 63368
rect 68100 63325 68109 63359
rect 68109 63325 68143 63359
rect 68143 63325 68152 63359
rect 68100 63316 68152 63325
rect 66444 63291 66496 63300
rect 66444 63257 66453 63291
rect 66453 63257 66487 63291
rect 66487 63257 66496 63291
rect 66444 63248 66496 63257
rect 19574 63078 19626 63130
rect 19638 63078 19690 63130
rect 19702 63078 19754 63130
rect 19766 63078 19818 63130
rect 19830 63078 19882 63130
rect 50294 63078 50346 63130
rect 50358 63078 50410 63130
rect 50422 63078 50474 63130
rect 50486 63078 50538 63130
rect 50550 63078 50602 63130
rect 23112 62883 23164 62892
rect 23112 62849 23121 62883
rect 23121 62849 23155 62883
rect 23155 62849 23164 62883
rect 23112 62840 23164 62849
rect 23388 62840 23440 62892
rect 24400 62840 24452 62892
rect 23848 62772 23900 62824
rect 56232 62976 56284 63028
rect 66444 62976 66496 63028
rect 24860 62908 24912 62960
rect 35348 62951 35400 62960
rect 35348 62917 35357 62951
rect 35357 62917 35391 62951
rect 35391 62917 35400 62951
rect 35348 62908 35400 62917
rect 35440 62908 35492 62960
rect 44180 62908 44232 62960
rect 36360 62840 36412 62892
rect 36452 62883 36504 62892
rect 36452 62849 36461 62883
rect 36461 62849 36495 62883
rect 36495 62849 36504 62883
rect 37648 62883 37700 62892
rect 36452 62840 36504 62849
rect 37648 62849 37657 62883
rect 37657 62849 37691 62883
rect 37691 62849 37700 62883
rect 37648 62840 37700 62849
rect 29092 62815 29144 62824
rect 29092 62781 29101 62815
rect 29101 62781 29135 62815
rect 29135 62781 29144 62815
rect 29092 62772 29144 62781
rect 29276 62772 29328 62824
rect 32956 62815 33008 62824
rect 32956 62781 32965 62815
rect 32965 62781 32999 62815
rect 32999 62781 33008 62815
rect 32956 62772 33008 62781
rect 33140 62815 33192 62824
rect 33140 62781 33149 62815
rect 33149 62781 33183 62815
rect 33183 62781 33192 62815
rect 33140 62772 33192 62781
rect 32496 62704 32548 62756
rect 35440 62636 35492 62688
rect 36084 62772 36136 62824
rect 36268 62815 36320 62824
rect 36268 62781 36277 62815
rect 36277 62781 36311 62815
rect 36311 62781 36320 62815
rect 36268 62772 36320 62781
rect 35716 62747 35768 62756
rect 35716 62713 35725 62747
rect 35725 62713 35759 62747
rect 35759 62713 35768 62747
rect 36636 62747 36688 62756
rect 35716 62704 35768 62713
rect 36636 62713 36645 62747
rect 36645 62713 36679 62747
rect 36679 62713 36688 62747
rect 36636 62704 36688 62713
rect 37924 62840 37976 62892
rect 57244 62840 57296 62892
rect 67548 62840 67600 62892
rect 38108 62772 38160 62824
rect 38016 62704 38068 62756
rect 35992 62636 36044 62688
rect 36176 62679 36228 62688
rect 36176 62645 36185 62679
rect 36185 62645 36219 62679
rect 36219 62645 36228 62679
rect 36176 62636 36228 62645
rect 38200 62636 38252 62688
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 34934 62534 34986 62586
rect 34998 62534 35050 62586
rect 35062 62534 35114 62586
rect 35126 62534 35178 62586
rect 35190 62534 35242 62586
rect 65654 62534 65706 62586
rect 65718 62534 65770 62586
rect 65782 62534 65834 62586
rect 65846 62534 65898 62586
rect 65910 62534 65962 62586
rect 23112 62432 23164 62484
rect 31024 62432 31076 62484
rect 33140 62475 33192 62484
rect 33140 62441 33149 62475
rect 33149 62441 33183 62475
rect 33183 62441 33192 62475
rect 33140 62432 33192 62441
rect 37924 62432 37976 62484
rect 35992 62364 36044 62416
rect 37648 62364 37700 62416
rect 23112 62339 23164 62348
rect 23112 62305 23121 62339
rect 23121 62305 23155 62339
rect 23155 62305 23164 62339
rect 23112 62296 23164 62305
rect 29368 62296 29420 62348
rect 21824 62228 21876 62280
rect 24400 62271 24452 62280
rect 24400 62237 24409 62271
rect 24409 62237 24443 62271
rect 24443 62237 24452 62271
rect 24400 62228 24452 62237
rect 26240 62271 26292 62280
rect 26240 62237 26249 62271
rect 26249 62237 26283 62271
rect 26283 62237 26292 62271
rect 26240 62228 26292 62237
rect 25320 62203 25372 62212
rect 25320 62169 25329 62203
rect 25329 62169 25363 62203
rect 25363 62169 25372 62203
rect 25320 62160 25372 62169
rect 25964 62160 26016 62212
rect 29000 62271 29052 62280
rect 29000 62237 29009 62271
rect 29009 62237 29043 62271
rect 29043 62237 29052 62271
rect 29000 62228 29052 62237
rect 29736 62271 29788 62280
rect 29736 62237 29745 62271
rect 29745 62237 29779 62271
rect 29779 62237 29788 62271
rect 29736 62228 29788 62237
rect 30380 62271 30432 62280
rect 30380 62237 30389 62271
rect 30389 62237 30423 62271
rect 30423 62237 30432 62271
rect 30380 62228 30432 62237
rect 26516 62203 26568 62212
rect 26516 62169 26550 62203
rect 26550 62169 26568 62203
rect 26516 62160 26568 62169
rect 19340 62092 19392 62144
rect 27436 62092 27488 62144
rect 28264 62135 28316 62144
rect 28264 62101 28273 62135
rect 28273 62101 28307 62135
rect 28307 62101 28316 62135
rect 28264 62092 28316 62101
rect 28816 62135 28868 62144
rect 28816 62101 28825 62135
rect 28825 62101 28859 62135
rect 28859 62101 28868 62135
rect 28816 62092 28868 62101
rect 29736 62092 29788 62144
rect 34704 62228 34756 62280
rect 35440 62296 35492 62348
rect 36636 62296 36688 62348
rect 35348 62271 35400 62280
rect 35348 62237 35357 62271
rect 35357 62237 35391 62271
rect 35391 62237 35400 62271
rect 38016 62271 38068 62280
rect 35348 62228 35400 62237
rect 38016 62237 38025 62271
rect 38025 62237 38059 62271
rect 38059 62237 38068 62271
rect 38016 62228 38068 62237
rect 38200 62271 38252 62280
rect 38200 62237 38209 62271
rect 38209 62237 38243 62271
rect 38243 62237 38252 62271
rect 38200 62228 38252 62237
rect 36636 62160 36688 62212
rect 66260 62228 66312 62280
rect 33692 62092 33744 62144
rect 35532 62135 35584 62144
rect 35532 62101 35541 62135
rect 35541 62101 35575 62135
rect 35575 62101 35584 62135
rect 35532 62092 35584 62101
rect 19574 61990 19626 62042
rect 19638 61990 19690 62042
rect 19702 61990 19754 62042
rect 19766 61990 19818 62042
rect 19830 61990 19882 62042
rect 50294 61990 50346 62042
rect 50358 61990 50410 62042
rect 50422 61990 50474 62042
rect 50486 61990 50538 62042
rect 50550 61990 50602 62042
rect 19340 61888 19392 61940
rect 26240 61888 26292 61940
rect 2964 61820 3016 61872
rect 25136 61863 25188 61872
rect 19340 61752 19392 61804
rect 20720 61752 20772 61804
rect 21824 61795 21876 61804
rect 21824 61761 21833 61795
rect 21833 61761 21867 61795
rect 21867 61761 21876 61795
rect 25136 61829 25145 61863
rect 25145 61829 25179 61863
rect 25179 61829 25188 61863
rect 25136 61820 25188 61829
rect 26056 61820 26108 61872
rect 21824 61752 21876 61761
rect 25688 61752 25740 61804
rect 25964 61795 26016 61804
rect 25964 61761 25973 61795
rect 25973 61761 26007 61795
rect 26007 61761 26016 61795
rect 25964 61752 26016 61761
rect 22744 61727 22796 61736
rect 22744 61693 22753 61727
rect 22753 61693 22787 61727
rect 22787 61693 22796 61727
rect 22744 61684 22796 61693
rect 23572 61684 23624 61736
rect 25872 61684 25924 61736
rect 38936 61888 38988 61940
rect 28816 61820 28868 61872
rect 28264 61752 28316 61804
rect 31760 61820 31812 61872
rect 30288 61752 30340 61804
rect 34796 61752 34848 61804
rect 33416 61727 33468 61736
rect 33416 61693 33425 61727
rect 33425 61693 33459 61727
rect 33459 61693 33468 61727
rect 33416 61684 33468 61693
rect 36452 61752 36504 61804
rect 66260 61820 66312 61872
rect 67640 61863 67692 61872
rect 67640 61829 67649 61863
rect 67649 61829 67683 61863
rect 67683 61829 67692 61863
rect 67640 61820 67692 61829
rect 35808 61727 35860 61736
rect 20352 61548 20404 61600
rect 21088 61591 21140 61600
rect 21088 61557 21097 61591
rect 21097 61557 21131 61591
rect 21131 61557 21140 61591
rect 21088 61548 21140 61557
rect 21180 61548 21232 61600
rect 24308 61548 24360 61600
rect 27804 61548 27856 61600
rect 27896 61548 27948 61600
rect 30380 61548 30432 61600
rect 34704 61548 34756 61600
rect 35808 61693 35817 61727
rect 35817 61693 35851 61727
rect 35851 61693 35860 61727
rect 35808 61684 35860 61693
rect 36084 61727 36136 61736
rect 36084 61693 36093 61727
rect 36093 61693 36127 61727
rect 36127 61693 36136 61727
rect 36084 61684 36136 61693
rect 35992 61616 36044 61668
rect 67640 61684 67692 61736
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 34934 61446 34986 61498
rect 34998 61446 35050 61498
rect 35062 61446 35114 61498
rect 35126 61446 35178 61498
rect 35190 61446 35242 61498
rect 65654 61446 65706 61498
rect 65718 61446 65770 61498
rect 65782 61446 65834 61498
rect 65846 61446 65898 61498
rect 65910 61446 65962 61498
rect 20352 61344 20404 61396
rect 20720 61387 20772 61396
rect 20720 61353 20729 61387
rect 20729 61353 20763 61387
rect 20763 61353 20772 61387
rect 20720 61344 20772 61353
rect 23572 61387 23624 61396
rect 23572 61353 23581 61387
rect 23581 61353 23615 61387
rect 23615 61353 23624 61387
rect 23572 61344 23624 61353
rect 26516 61344 26568 61396
rect 29000 61344 29052 61396
rect 19616 61276 19668 61328
rect 19432 61251 19484 61260
rect 19432 61217 19441 61251
rect 19441 61217 19475 61251
rect 19475 61217 19484 61251
rect 19432 61208 19484 61217
rect 18236 61140 18288 61192
rect 19616 61183 19668 61192
rect 19616 61149 19625 61183
rect 19625 61149 19659 61183
rect 19659 61149 19668 61183
rect 19616 61140 19668 61149
rect 19984 61004 20036 61056
rect 27804 61276 27856 61328
rect 29736 61276 29788 61328
rect 21180 61251 21232 61260
rect 21180 61217 21189 61251
rect 21189 61217 21223 61251
rect 21223 61217 21232 61251
rect 21180 61208 21232 61217
rect 21088 61140 21140 61192
rect 24860 61208 24912 61260
rect 24400 61183 24452 61192
rect 24400 61149 24409 61183
rect 24409 61149 24443 61183
rect 24443 61149 24452 61183
rect 24400 61140 24452 61149
rect 27436 61183 27488 61192
rect 27436 61149 27445 61183
rect 27445 61149 27479 61183
rect 27479 61149 27488 61183
rect 27436 61140 27488 61149
rect 25872 61072 25924 61124
rect 27896 61140 27948 61192
rect 28356 61140 28408 61192
rect 32956 61344 33008 61396
rect 33416 61344 33468 61396
rect 67640 61387 67692 61396
rect 34796 61319 34848 61328
rect 34796 61285 34805 61319
rect 34805 61285 34839 61319
rect 34839 61285 34848 61319
rect 34796 61276 34848 61285
rect 36084 61276 36136 61328
rect 31484 61208 31536 61260
rect 31024 61183 31076 61192
rect 31024 61149 31033 61183
rect 31033 61149 31067 61183
rect 31067 61149 31076 61183
rect 31024 61140 31076 61149
rect 31208 61183 31260 61192
rect 31208 61149 31217 61183
rect 31217 61149 31251 61183
rect 31251 61149 31260 61183
rect 31208 61140 31260 61149
rect 31760 61140 31812 61192
rect 32404 61140 32456 61192
rect 34704 61140 34756 61192
rect 35072 61183 35124 61192
rect 35072 61149 35081 61183
rect 35081 61149 35115 61183
rect 35115 61149 35124 61183
rect 35072 61140 35124 61149
rect 35348 61140 35400 61192
rect 35992 61183 36044 61192
rect 35992 61149 36001 61183
rect 36001 61149 36035 61183
rect 36035 61149 36044 61183
rect 35992 61140 36044 61149
rect 36176 61183 36228 61192
rect 36176 61149 36185 61183
rect 36185 61149 36219 61183
rect 36219 61149 36228 61183
rect 36360 61183 36412 61192
rect 36176 61140 36228 61149
rect 36360 61149 36369 61183
rect 36369 61149 36403 61183
rect 36403 61149 36412 61183
rect 36360 61140 36412 61149
rect 67640 61353 67649 61387
rect 67649 61353 67683 61387
rect 67683 61353 67692 61387
rect 67640 61344 67692 61353
rect 37372 61140 37424 61192
rect 38108 61140 38160 61192
rect 39948 61140 40000 61192
rect 67548 61183 67600 61192
rect 67548 61149 67557 61183
rect 67557 61149 67591 61183
rect 67591 61149 67600 61183
rect 67548 61140 67600 61149
rect 35532 61072 35584 61124
rect 20812 61004 20864 61056
rect 38752 61115 38804 61124
rect 38752 61081 38761 61115
rect 38761 61081 38795 61115
rect 38795 61081 38804 61115
rect 38752 61072 38804 61081
rect 40132 61115 40184 61124
rect 40132 61081 40166 61115
rect 40166 61081 40184 61115
rect 40132 61072 40184 61081
rect 36544 61004 36596 61056
rect 41236 61047 41288 61056
rect 41236 61013 41245 61047
rect 41245 61013 41279 61047
rect 41279 61013 41288 61047
rect 41236 61004 41288 61013
rect 19574 60902 19626 60954
rect 19638 60902 19690 60954
rect 19702 60902 19754 60954
rect 19766 60902 19818 60954
rect 19830 60902 19882 60954
rect 50294 60902 50346 60954
rect 50358 60902 50410 60954
rect 50422 60902 50474 60954
rect 50486 60902 50538 60954
rect 50550 60902 50602 60954
rect 19340 60800 19392 60852
rect 26240 60843 26292 60852
rect 26240 60809 26249 60843
rect 26249 60809 26283 60843
rect 26283 60809 26292 60843
rect 30288 60843 30340 60852
rect 26240 60800 26292 60809
rect 30288 60809 30297 60843
rect 30297 60809 30331 60843
rect 30331 60809 30340 60843
rect 30288 60800 30340 60809
rect 36360 60800 36412 60852
rect 40132 60800 40184 60852
rect 1860 60775 1912 60784
rect 1860 60741 1869 60775
rect 1869 60741 1903 60775
rect 1903 60741 1912 60775
rect 1860 60732 1912 60741
rect 17040 60664 17092 60716
rect 17500 60664 17552 60716
rect 19984 60664 20036 60716
rect 17408 60639 17460 60648
rect 17408 60605 17417 60639
rect 17417 60605 17451 60639
rect 17451 60605 17460 60639
rect 17408 60596 17460 60605
rect 22008 60596 22060 60648
rect 25504 60664 25556 60716
rect 26332 60596 26384 60648
rect 27712 60664 27764 60716
rect 30380 60664 30432 60716
rect 31484 60732 31536 60784
rect 2136 60503 2188 60512
rect 2136 60469 2145 60503
rect 2145 60469 2179 60503
rect 2179 60469 2188 60503
rect 2136 60460 2188 60469
rect 15844 60460 15896 60512
rect 16028 60460 16080 60512
rect 23664 60528 23716 60580
rect 30472 60596 30524 60648
rect 18788 60503 18840 60512
rect 18788 60469 18797 60503
rect 18797 60469 18831 60503
rect 18831 60469 18840 60503
rect 18788 60460 18840 60469
rect 21548 60460 21600 60512
rect 22376 60460 22428 60512
rect 22836 60460 22888 60512
rect 24952 60503 25004 60512
rect 24952 60469 24961 60503
rect 24961 60469 24995 60503
rect 24995 60469 25004 60503
rect 24952 60460 25004 60469
rect 28080 60528 28132 60580
rect 31208 60664 31260 60716
rect 33692 60707 33744 60716
rect 33692 60673 33701 60707
rect 33701 60673 33735 60707
rect 33735 60673 33744 60707
rect 33692 60664 33744 60673
rect 36084 60664 36136 60716
rect 36544 60707 36596 60716
rect 36544 60673 36553 60707
rect 36553 60673 36587 60707
rect 36587 60673 36596 60707
rect 36544 60664 36596 60673
rect 38108 60707 38160 60716
rect 35992 60596 36044 60648
rect 38108 60673 38117 60707
rect 38117 60673 38151 60707
rect 38151 60673 38160 60707
rect 38108 60664 38160 60673
rect 38660 60664 38712 60716
rect 39856 60664 39908 60716
rect 40132 60707 40184 60716
rect 40132 60673 40141 60707
rect 40141 60673 40175 60707
rect 40175 60673 40184 60707
rect 40132 60664 40184 60673
rect 35072 60528 35124 60580
rect 67364 60596 67416 60648
rect 67548 60639 67600 60648
rect 67548 60605 67557 60639
rect 67557 60605 67591 60639
rect 67591 60605 67600 60639
rect 67548 60596 67600 60605
rect 68100 60528 68152 60580
rect 33968 60460 34020 60512
rect 39212 60460 39264 60512
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 65654 60358 65706 60410
rect 65718 60358 65770 60410
rect 65782 60358 65834 60410
rect 65846 60358 65898 60410
rect 65910 60358 65962 60410
rect 19984 60256 20036 60308
rect 19248 60188 19300 60240
rect 18788 60120 18840 60172
rect 20812 60163 20864 60172
rect 20812 60129 20821 60163
rect 20821 60129 20855 60163
rect 20855 60129 20864 60163
rect 20812 60120 20864 60129
rect 21548 60120 21600 60172
rect 25780 60299 25832 60308
rect 25780 60265 25789 60299
rect 25789 60265 25823 60299
rect 25823 60265 25832 60299
rect 25780 60256 25832 60265
rect 28264 60256 28316 60308
rect 30472 60256 30524 60308
rect 31024 60256 31076 60308
rect 38660 60256 38712 60308
rect 40132 60256 40184 60308
rect 67364 60299 67416 60308
rect 67364 60265 67373 60299
rect 67373 60265 67407 60299
rect 67407 60265 67416 60299
rect 67364 60256 67416 60265
rect 68100 60299 68152 60308
rect 68100 60265 68109 60299
rect 68109 60265 68143 60299
rect 68143 60265 68152 60299
rect 68100 60256 68152 60265
rect 27620 60188 27672 60240
rect 27436 60120 27488 60172
rect 27804 60163 27856 60172
rect 27804 60129 27813 60163
rect 27813 60129 27847 60163
rect 27847 60129 27856 60163
rect 27804 60120 27856 60129
rect 28264 60120 28316 60172
rect 1676 60052 1728 60104
rect 15568 60095 15620 60104
rect 15568 60061 15577 60095
rect 15577 60061 15611 60095
rect 15611 60061 15620 60095
rect 15568 60052 15620 60061
rect 15844 60095 15896 60104
rect 15844 60061 15878 60095
rect 15878 60061 15896 60095
rect 15844 60052 15896 60061
rect 16580 60052 16632 60104
rect 20996 60095 21048 60104
rect 20996 60061 21005 60095
rect 21005 60061 21039 60095
rect 21039 60061 21048 60095
rect 20996 60052 21048 60061
rect 21732 60095 21784 60104
rect 21732 60061 21741 60095
rect 21741 60061 21775 60095
rect 21775 60061 21784 60095
rect 23756 60095 23808 60104
rect 21732 60052 21784 60061
rect 23756 60061 23765 60095
rect 23765 60061 23799 60095
rect 23799 60061 23808 60095
rect 23756 60052 23808 60061
rect 24952 60052 25004 60104
rect 26332 60095 26384 60104
rect 26332 60061 26341 60095
rect 26341 60061 26375 60095
rect 26375 60061 26384 60095
rect 26332 60052 26384 60061
rect 16948 59959 17000 59968
rect 16948 59925 16957 59959
rect 16957 59925 16991 59959
rect 16991 59925 17000 59959
rect 16948 59916 17000 59925
rect 17592 59916 17644 59968
rect 17868 59916 17920 59968
rect 26332 59916 26384 59968
rect 26976 59916 27028 59968
rect 28080 60095 28132 60104
rect 28080 60061 28089 60095
rect 28089 60061 28123 60095
rect 28123 60061 28132 60095
rect 28540 60120 28592 60172
rect 28080 60052 28132 60061
rect 29920 60052 29972 60104
rect 38844 60120 38896 60172
rect 39948 60120 40000 60172
rect 31668 60052 31720 60104
rect 31760 60095 31812 60104
rect 31760 60061 31769 60095
rect 31769 60061 31803 60095
rect 31803 60061 31812 60095
rect 31760 60052 31812 60061
rect 32404 60052 32456 60104
rect 36544 60052 36596 60104
rect 38936 60095 38988 60104
rect 38936 60061 38945 60095
rect 38945 60061 38979 60095
rect 38979 60061 38988 60095
rect 38936 60052 38988 60061
rect 39672 60052 39724 60104
rect 40132 60095 40184 60104
rect 40132 60061 40141 60095
rect 40141 60061 40175 60095
rect 40175 60061 40184 60095
rect 40132 60052 40184 60061
rect 42708 60052 42760 60104
rect 32220 59984 32272 60036
rect 33048 59984 33100 60036
rect 40224 59984 40276 60036
rect 41236 59984 41288 60036
rect 44088 59984 44140 60036
rect 29276 59916 29328 59968
rect 29644 59916 29696 59968
rect 31852 59916 31904 59968
rect 33784 59916 33836 59968
rect 35348 59959 35400 59968
rect 35348 59925 35357 59959
rect 35357 59925 35391 59959
rect 35391 59925 35400 59959
rect 35348 59916 35400 59925
rect 42984 59916 43036 59968
rect 19574 59814 19626 59866
rect 19638 59814 19690 59866
rect 19702 59814 19754 59866
rect 19766 59814 19818 59866
rect 19830 59814 19882 59866
rect 50294 59814 50346 59866
rect 50358 59814 50410 59866
rect 50422 59814 50474 59866
rect 50486 59814 50538 59866
rect 50550 59814 50602 59866
rect 15568 59712 15620 59764
rect 17040 59755 17092 59764
rect 17040 59721 17049 59755
rect 17049 59721 17083 59755
rect 17083 59721 17092 59755
rect 17040 59712 17092 59721
rect 17408 59712 17460 59764
rect 1676 59619 1728 59628
rect 1676 59585 1685 59619
rect 1685 59585 1719 59619
rect 1719 59585 1728 59619
rect 1676 59576 1728 59585
rect 14648 59619 14700 59628
rect 14648 59585 14657 59619
rect 14657 59585 14691 59619
rect 14691 59585 14700 59619
rect 14648 59576 14700 59585
rect 15844 59619 15896 59628
rect 15844 59585 15853 59619
rect 15853 59585 15887 59619
rect 15887 59585 15896 59619
rect 15844 59576 15896 59585
rect 16580 59576 16632 59628
rect 17868 59576 17920 59628
rect 19432 59712 19484 59764
rect 25504 59755 25556 59764
rect 25504 59721 25513 59755
rect 25513 59721 25547 59755
rect 25547 59721 25556 59755
rect 25504 59712 25556 59721
rect 26332 59712 26384 59764
rect 18788 59619 18840 59628
rect 18788 59585 18797 59619
rect 18797 59585 18831 59619
rect 18831 59585 18840 59619
rect 18788 59576 18840 59585
rect 19524 59619 19576 59628
rect 19524 59585 19533 59619
rect 19533 59585 19567 59619
rect 19567 59585 19576 59619
rect 22376 59619 22428 59628
rect 19524 59576 19576 59585
rect 22376 59585 22385 59619
rect 22385 59585 22419 59619
rect 22419 59585 22428 59619
rect 22376 59576 22428 59585
rect 22836 59619 22888 59628
rect 22836 59585 22845 59619
rect 22845 59585 22879 59619
rect 22879 59585 22888 59619
rect 22836 59576 22888 59585
rect 25780 59644 25832 59696
rect 26240 59644 26292 59696
rect 28080 59712 28132 59764
rect 32220 59755 32272 59764
rect 32220 59721 32229 59755
rect 32229 59721 32263 59755
rect 32263 59721 32272 59755
rect 32220 59712 32272 59721
rect 36544 59755 36596 59764
rect 36544 59721 36553 59755
rect 36553 59721 36587 59755
rect 36587 59721 36596 59755
rect 36544 59712 36596 59721
rect 44088 59755 44140 59764
rect 44088 59721 44097 59755
rect 44097 59721 44131 59755
rect 44131 59721 44140 59755
rect 44088 59712 44140 59721
rect 31760 59644 31812 59696
rect 33968 59687 34020 59696
rect 25412 59576 25464 59628
rect 26976 59619 27028 59628
rect 26976 59585 26985 59619
rect 26985 59585 27019 59619
rect 27019 59585 27028 59619
rect 26976 59576 27028 59585
rect 27620 59576 27672 59628
rect 28540 59576 28592 59628
rect 28908 59576 28960 59628
rect 29644 59619 29696 59628
rect 29644 59585 29678 59619
rect 29678 59585 29696 59619
rect 29644 59576 29696 59585
rect 33968 59653 33977 59687
rect 33977 59653 34011 59687
rect 34011 59653 34020 59687
rect 33968 59644 34020 59653
rect 53840 59644 53892 59696
rect 1860 59551 1912 59560
rect 1860 59517 1869 59551
rect 1869 59517 1903 59551
rect 1903 59517 1912 59551
rect 1860 59508 1912 59517
rect 2780 59551 2832 59560
rect 2780 59517 2789 59551
rect 2789 59517 2823 59551
rect 2823 59517 2832 59551
rect 2780 59508 2832 59517
rect 16948 59508 17000 59560
rect 19984 59508 20036 59560
rect 29368 59551 29420 59560
rect 29368 59517 29377 59551
rect 29377 59517 29411 59551
rect 29411 59517 29420 59551
rect 29368 59508 29420 59517
rect 31576 59508 31628 59560
rect 32680 59619 32732 59628
rect 32680 59585 32689 59619
rect 32689 59585 32723 59619
rect 32723 59585 32732 59619
rect 32680 59576 32732 59585
rect 32864 59619 32916 59628
rect 32864 59585 32873 59619
rect 32873 59585 32907 59619
rect 32907 59585 32916 59619
rect 33784 59619 33836 59628
rect 32864 59576 32916 59585
rect 33784 59585 33793 59619
rect 33793 59585 33827 59619
rect 33827 59585 33836 59619
rect 33784 59576 33836 59585
rect 37372 59576 37424 59628
rect 39672 59619 39724 59628
rect 39672 59585 39681 59619
rect 39681 59585 39715 59619
rect 39715 59585 39724 59619
rect 39672 59576 39724 59585
rect 41604 59619 41656 59628
rect 35992 59508 36044 59560
rect 36268 59508 36320 59560
rect 37280 59551 37332 59560
rect 37280 59517 37289 59551
rect 37289 59517 37323 59551
rect 37323 59517 37332 59551
rect 37280 59508 37332 59517
rect 39212 59508 39264 59560
rect 41604 59585 41613 59619
rect 41613 59585 41647 59619
rect 41647 59585 41656 59619
rect 41604 59576 41656 59585
rect 41696 59619 41748 59628
rect 41696 59585 41705 59619
rect 41705 59585 41739 59619
rect 41739 59585 41748 59619
rect 41696 59576 41748 59585
rect 42984 59576 43036 59628
rect 43536 59576 43588 59628
rect 44180 59619 44232 59628
rect 44180 59585 44189 59619
rect 44189 59585 44223 59619
rect 44223 59585 44232 59619
rect 44180 59576 44232 59585
rect 67272 59619 67324 59628
rect 67272 59585 67281 59619
rect 67281 59585 67315 59619
rect 67315 59585 67324 59619
rect 67272 59576 67324 59585
rect 41512 59508 41564 59560
rect 42616 59508 42668 59560
rect 19248 59483 19300 59492
rect 19248 59449 19257 59483
rect 19257 59449 19291 59483
rect 19291 59449 19300 59483
rect 19248 59440 19300 59449
rect 22192 59440 22244 59492
rect 36360 59483 36412 59492
rect 36360 59449 36369 59483
rect 36369 59449 36403 59483
rect 36403 59449 36412 59483
rect 36360 59440 36412 59449
rect 36636 59440 36688 59492
rect 42708 59440 42760 59492
rect 14372 59372 14424 59424
rect 18788 59372 18840 59424
rect 20352 59372 20404 59424
rect 22008 59372 22060 59424
rect 29276 59372 29328 59424
rect 39120 59372 39172 59424
rect 41420 59415 41472 59424
rect 41420 59381 41429 59415
rect 41429 59381 41463 59415
rect 41463 59381 41472 59415
rect 41420 59372 41472 59381
rect 43076 59372 43128 59424
rect 43168 59372 43220 59424
rect 67180 59372 67232 59424
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 34934 59270 34986 59322
rect 34998 59270 35050 59322
rect 35062 59270 35114 59322
rect 35126 59270 35178 59322
rect 35190 59270 35242 59322
rect 65654 59270 65706 59322
rect 65718 59270 65770 59322
rect 65782 59270 65834 59322
rect 65846 59270 65898 59322
rect 65910 59270 65962 59322
rect 1860 59168 1912 59220
rect 17500 59168 17552 59220
rect 15476 59143 15528 59152
rect 15476 59109 15485 59143
rect 15485 59109 15519 59143
rect 15519 59109 15528 59143
rect 15476 59100 15528 59109
rect 19524 59100 19576 59152
rect 2044 58964 2096 59016
rect 6000 58964 6052 59016
rect 14096 59007 14148 59016
rect 14096 58973 14105 59007
rect 14105 58973 14139 59007
rect 14139 58973 14148 59007
rect 14096 58964 14148 58973
rect 14372 59007 14424 59016
rect 14372 58973 14406 59007
rect 14406 58973 14424 59007
rect 14372 58964 14424 58973
rect 17592 59007 17644 59016
rect 17592 58973 17601 59007
rect 17601 58973 17635 59007
rect 17635 58973 17644 59007
rect 17592 58964 17644 58973
rect 19432 59007 19484 59016
rect 19432 58973 19441 59007
rect 19441 58973 19475 59007
rect 19475 58973 19484 59007
rect 19432 58964 19484 58973
rect 20168 59007 20220 59016
rect 20168 58973 20177 59007
rect 20177 58973 20211 59007
rect 20211 58973 20220 59007
rect 20168 58964 20220 58973
rect 21272 58964 21324 59016
rect 20444 58896 20496 58948
rect 29920 59211 29972 59220
rect 29920 59177 29929 59211
rect 29929 59177 29963 59211
rect 29963 59177 29972 59211
rect 29920 59168 29972 59177
rect 32680 59168 32732 59220
rect 36268 59211 36320 59220
rect 36268 59177 36277 59211
rect 36277 59177 36311 59211
rect 36311 59177 36320 59211
rect 36268 59168 36320 59177
rect 39856 59211 39908 59220
rect 39856 59177 39865 59211
rect 39865 59177 39899 59211
rect 39899 59177 39908 59211
rect 39856 59168 39908 59177
rect 41604 59168 41656 59220
rect 25596 58964 25648 59016
rect 31668 59007 31720 59016
rect 31668 58973 31677 59007
rect 31677 58973 31711 59007
rect 31711 58973 31720 59007
rect 31668 58964 31720 58973
rect 37280 59032 37332 59084
rect 39120 59075 39172 59084
rect 39120 59041 39129 59075
rect 39129 59041 39163 59075
rect 39163 59041 39172 59075
rect 39120 59032 39172 59041
rect 39672 59032 39724 59084
rect 40224 59075 40276 59084
rect 40224 59041 40233 59075
rect 40233 59041 40267 59075
rect 40267 59041 40276 59075
rect 40224 59032 40276 59041
rect 38844 59007 38896 59016
rect 29276 58896 29328 58948
rect 30932 58896 30984 58948
rect 35348 58896 35400 58948
rect 38844 58973 38853 59007
rect 38853 58973 38887 59007
rect 38887 58973 38896 59007
rect 38844 58964 38896 58973
rect 38016 58896 38068 58948
rect 39948 58964 40000 59016
rect 40316 59007 40368 59016
rect 40316 58973 40325 59007
rect 40325 58973 40359 59007
rect 40359 58973 40368 59007
rect 40316 58964 40368 58973
rect 40776 58964 40828 59016
rect 44180 59168 44232 59220
rect 42616 59032 42668 59084
rect 42708 58964 42760 59016
rect 43444 58964 43496 59016
rect 40224 58896 40276 58948
rect 41236 58896 41288 58948
rect 42984 58939 43036 58948
rect 42984 58905 42993 58939
rect 42993 58905 43027 58939
rect 43027 58905 43036 58939
rect 42984 58896 43036 58905
rect 19064 58828 19116 58880
rect 19984 58871 20036 58880
rect 19984 58837 19993 58871
rect 19993 58837 20027 58871
rect 20027 58837 20036 58871
rect 19984 58828 20036 58837
rect 21456 58871 21508 58880
rect 21456 58837 21465 58871
rect 21465 58837 21499 58871
rect 21499 58837 21508 58871
rect 21456 58828 21508 58837
rect 25228 58871 25280 58880
rect 25228 58837 25237 58871
rect 25237 58837 25271 58871
rect 25271 58837 25280 58871
rect 25228 58828 25280 58837
rect 30472 58828 30524 58880
rect 31760 58828 31812 58880
rect 37464 58828 37516 58880
rect 38844 58828 38896 58880
rect 39948 58828 40000 58880
rect 19574 58726 19626 58778
rect 19638 58726 19690 58778
rect 19702 58726 19754 58778
rect 19766 58726 19818 58778
rect 19830 58726 19882 58778
rect 50294 58726 50346 58778
rect 50358 58726 50410 58778
rect 50422 58726 50474 58778
rect 50486 58726 50538 58778
rect 50550 58726 50602 58778
rect 14096 58667 14148 58676
rect 14096 58633 14105 58667
rect 14105 58633 14139 58667
rect 14139 58633 14148 58667
rect 14096 58624 14148 58633
rect 14648 58624 14700 58676
rect 20352 58624 20404 58676
rect 20628 58624 20680 58676
rect 21272 58667 21324 58676
rect 21272 58633 21281 58667
rect 21281 58633 21315 58667
rect 21315 58633 21324 58667
rect 21272 58624 21324 58633
rect 13820 58488 13872 58540
rect 15476 58556 15528 58608
rect 19984 58556 20036 58608
rect 20996 58556 21048 58608
rect 15200 58488 15252 58540
rect 16028 58488 16080 58540
rect 17132 58531 17184 58540
rect 17132 58497 17141 58531
rect 17141 58497 17175 58531
rect 17175 58497 17184 58531
rect 17132 58488 17184 58497
rect 19064 58531 19116 58540
rect 19064 58497 19073 58531
rect 19073 58497 19107 58531
rect 19107 58497 19116 58531
rect 19064 58488 19116 58497
rect 25596 58667 25648 58676
rect 25596 58633 25605 58667
rect 25605 58633 25639 58667
rect 25639 58633 25648 58667
rect 25596 58624 25648 58633
rect 26240 58624 26292 58676
rect 28908 58624 28960 58676
rect 31760 58624 31812 58676
rect 37372 58624 37424 58676
rect 39672 58624 39724 58676
rect 41236 58667 41288 58676
rect 41236 58633 41245 58667
rect 41245 58633 41279 58667
rect 41279 58633 41288 58667
rect 41236 58624 41288 58633
rect 21456 58556 21508 58608
rect 24308 58531 24360 58540
rect 24308 58497 24317 58531
rect 24317 58497 24351 58531
rect 24351 58497 24360 58531
rect 24308 58488 24360 58497
rect 27804 58556 27856 58608
rect 25412 58531 25464 58540
rect 25412 58497 25421 58531
rect 25421 58497 25455 58531
rect 25455 58497 25464 58531
rect 25412 58488 25464 58497
rect 26424 58488 26476 58540
rect 27712 58488 27764 58540
rect 27896 58531 27948 58540
rect 27896 58497 27905 58531
rect 27905 58497 27939 58531
rect 27939 58497 27948 58531
rect 27896 58488 27948 58497
rect 20996 58420 21048 58472
rect 28908 58531 28960 58540
rect 28908 58497 28942 58531
rect 28942 58497 28960 58531
rect 29092 58531 29144 58540
rect 28908 58488 28960 58497
rect 29092 58497 29101 58531
rect 29101 58497 29135 58531
rect 29135 58497 29144 58531
rect 29092 58488 29144 58497
rect 29828 58488 29880 58540
rect 31300 58531 31352 58540
rect 31300 58497 31309 58531
rect 31309 58497 31343 58531
rect 31343 58497 31352 58531
rect 31300 58488 31352 58497
rect 31668 58488 31720 58540
rect 35348 58556 35400 58608
rect 38752 58556 38804 58608
rect 33692 58488 33744 58540
rect 37464 58531 37516 58540
rect 37464 58497 37473 58531
rect 37473 58497 37507 58531
rect 37507 58497 37516 58531
rect 37464 58488 37516 58497
rect 39120 58556 39172 58608
rect 41512 58556 41564 58608
rect 39212 58531 39264 58540
rect 39212 58497 39221 58531
rect 39221 58497 39255 58531
rect 39255 58497 39264 58531
rect 39212 58488 39264 58497
rect 39948 58488 40000 58540
rect 40316 58488 40368 58540
rect 28540 58463 28592 58472
rect 16764 58284 16816 58336
rect 20444 58284 20496 58336
rect 24584 58284 24636 58336
rect 26332 58327 26384 58336
rect 26332 58293 26341 58327
rect 26341 58293 26375 58327
rect 26375 58293 26384 58327
rect 26332 58284 26384 58293
rect 26976 58284 27028 58336
rect 28540 58429 28549 58463
rect 28549 58429 28583 58463
rect 28583 58429 28592 58463
rect 28540 58420 28592 58429
rect 28816 58463 28868 58472
rect 28816 58429 28825 58463
rect 28825 58429 28859 58463
rect 28859 58429 28868 58463
rect 28816 58420 28868 58429
rect 40224 58420 40276 58472
rect 41420 58531 41472 58540
rect 41420 58497 41429 58531
rect 41429 58497 41463 58531
rect 41463 58497 41472 58531
rect 41420 58488 41472 58497
rect 41604 58488 41656 58540
rect 42984 58488 43036 58540
rect 43168 58420 43220 58472
rect 43444 58463 43496 58472
rect 43444 58429 43453 58463
rect 43453 58429 43487 58463
rect 43487 58429 43496 58463
rect 43444 58420 43496 58429
rect 38936 58352 38988 58404
rect 42708 58352 42760 58404
rect 43720 58463 43772 58472
rect 43720 58429 43729 58463
rect 43729 58429 43763 58463
rect 43763 58429 43772 58463
rect 43720 58420 43772 58429
rect 43904 58420 43956 58472
rect 29920 58284 29972 58336
rect 30380 58327 30432 58336
rect 30380 58293 30389 58327
rect 30389 58293 30423 58327
rect 30423 58293 30432 58327
rect 30380 58284 30432 58293
rect 31116 58327 31168 58336
rect 31116 58293 31125 58327
rect 31125 58293 31159 58327
rect 31159 58293 31168 58327
rect 31116 58284 31168 58293
rect 32588 58284 32640 58336
rect 33876 58284 33928 58336
rect 38660 58284 38712 58336
rect 41420 58284 41472 58336
rect 41604 58327 41656 58336
rect 41604 58293 41613 58327
rect 41613 58293 41647 58327
rect 41647 58293 41656 58327
rect 41604 58284 41656 58293
rect 44272 58284 44324 58336
rect 66260 58284 66312 58336
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 34934 58182 34986 58234
rect 34998 58182 35050 58234
rect 35062 58182 35114 58234
rect 35126 58182 35178 58234
rect 35190 58182 35242 58234
rect 65654 58182 65706 58234
rect 65718 58182 65770 58234
rect 65782 58182 65834 58234
rect 65846 58182 65898 58234
rect 65910 58182 65962 58234
rect 20168 58123 20220 58132
rect 20168 58089 20177 58123
rect 20177 58089 20211 58123
rect 20211 58089 20220 58123
rect 20168 58080 20220 58089
rect 20996 58123 21048 58132
rect 20996 58089 21005 58123
rect 21005 58089 21039 58123
rect 21039 58089 21048 58123
rect 20996 58080 21048 58089
rect 28080 58123 28132 58132
rect 28080 58089 28089 58123
rect 28089 58089 28123 58123
rect 28123 58089 28132 58123
rect 28080 58080 28132 58089
rect 28816 58080 28868 58132
rect 38016 58080 38068 58132
rect 43904 58080 43956 58132
rect 20444 58012 20496 58064
rect 39028 58012 39080 58064
rect 24584 57987 24636 57996
rect 24584 57953 24593 57987
rect 24593 57953 24627 57987
rect 24627 57953 24636 57987
rect 24584 57944 24636 57953
rect 26148 57987 26200 57996
rect 26148 57953 26157 57987
rect 26157 57953 26191 57987
rect 26191 57953 26200 57987
rect 26148 57944 26200 57953
rect 26332 57944 26384 57996
rect 15844 57919 15896 57928
rect 15844 57885 15853 57919
rect 15853 57885 15887 57919
rect 15887 57885 15896 57919
rect 15844 57876 15896 57885
rect 16764 57919 16816 57928
rect 16764 57885 16798 57919
rect 16798 57885 16816 57919
rect 16764 57876 16816 57885
rect 19432 57876 19484 57928
rect 22468 57919 22520 57928
rect 22468 57885 22477 57919
rect 22477 57885 22511 57919
rect 22511 57885 22520 57919
rect 22468 57876 22520 57885
rect 20352 57808 20404 57860
rect 22744 57851 22796 57860
rect 22744 57817 22778 57851
rect 22778 57817 22796 57851
rect 22744 57808 22796 57817
rect 17868 57783 17920 57792
rect 17868 57749 17877 57783
rect 17877 57749 17911 57783
rect 17911 57749 17920 57783
rect 17868 57740 17920 57749
rect 19156 57740 19208 57792
rect 19984 57783 20036 57792
rect 19984 57749 20009 57783
rect 20009 57749 20036 57783
rect 19984 57740 20036 57749
rect 20628 57740 20680 57792
rect 23020 57740 23072 57792
rect 26976 57919 27028 57928
rect 26976 57885 27010 57919
rect 27010 57885 27028 57919
rect 26976 57876 27028 57885
rect 29828 57876 29880 57928
rect 30380 57876 30432 57928
rect 31116 57876 31168 57928
rect 33048 57876 33100 57928
rect 36268 57876 36320 57928
rect 37648 57876 37700 57928
rect 38660 57876 38712 57928
rect 38844 57876 38896 57928
rect 44272 57919 44324 57928
rect 44272 57885 44281 57919
rect 44281 57885 44315 57919
rect 44315 57885 44324 57919
rect 44272 57876 44324 57885
rect 66260 57919 66312 57928
rect 29368 57808 29420 57860
rect 32128 57808 32180 57860
rect 33968 57808 34020 57860
rect 43076 57808 43128 57860
rect 66260 57885 66269 57919
rect 66269 57885 66303 57919
rect 66303 57885 66312 57919
rect 66260 57876 66312 57885
rect 68100 57919 68152 57928
rect 68100 57885 68109 57919
rect 68109 57885 68143 57919
rect 68143 57885 68152 57919
rect 68100 57876 68152 57885
rect 29920 57740 29972 57792
rect 33692 57740 33744 57792
rect 36084 57783 36136 57792
rect 36084 57749 36093 57783
rect 36093 57749 36127 57783
rect 36127 57749 36136 57783
rect 36084 57740 36136 57749
rect 36544 57740 36596 57792
rect 66444 57851 66496 57860
rect 66444 57817 66453 57851
rect 66453 57817 66487 57851
rect 66487 57817 66496 57851
rect 66444 57808 66496 57817
rect 46388 57783 46440 57792
rect 46388 57749 46397 57783
rect 46397 57749 46431 57783
rect 46431 57749 46440 57783
rect 46388 57740 46440 57749
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 17132 57536 17184 57588
rect 14924 57400 14976 57452
rect 17868 57468 17920 57520
rect 19340 57536 19392 57588
rect 22468 57536 22520 57588
rect 33048 57536 33100 57588
rect 36268 57536 36320 57588
rect 37556 57536 37608 57588
rect 40776 57536 40828 57588
rect 66444 57536 66496 57588
rect 22744 57511 22796 57520
rect 22744 57477 22753 57511
rect 22753 57477 22787 57511
rect 22787 57477 22796 57511
rect 22744 57468 22796 57477
rect 25228 57468 25280 57520
rect 27712 57468 27764 57520
rect 29920 57511 29972 57520
rect 29920 57477 29929 57511
rect 29929 57477 29963 57511
rect 29963 57477 29972 57511
rect 29920 57468 29972 57477
rect 30472 57468 30524 57520
rect 32128 57511 32180 57520
rect 32128 57477 32137 57511
rect 32137 57477 32171 57511
rect 32171 57477 32180 57511
rect 32128 57468 32180 57477
rect 33876 57511 33928 57520
rect 14372 57375 14424 57384
rect 14372 57341 14381 57375
rect 14381 57341 14415 57375
rect 14415 57341 14424 57375
rect 14372 57332 14424 57341
rect 16580 57332 16632 57384
rect 19156 57443 19208 57452
rect 19156 57409 19190 57443
rect 19190 57409 19208 57443
rect 23020 57443 23072 57452
rect 19156 57400 19208 57409
rect 23020 57409 23029 57443
rect 23029 57409 23063 57443
rect 23063 57409 23072 57443
rect 23020 57400 23072 57409
rect 18144 57375 18196 57384
rect 18144 57341 18153 57375
rect 18153 57341 18187 57375
rect 18187 57341 18196 57375
rect 18144 57332 18196 57341
rect 15752 57307 15804 57316
rect 15752 57273 15761 57307
rect 15761 57273 15795 57307
rect 15795 57273 15804 57307
rect 20076 57332 20128 57384
rect 23204 57443 23256 57452
rect 23204 57409 23213 57443
rect 23213 57409 23247 57443
rect 23247 57409 23256 57443
rect 23204 57400 23256 57409
rect 23664 57400 23716 57452
rect 24952 57400 25004 57452
rect 27620 57443 27672 57452
rect 27620 57409 27629 57443
rect 27629 57409 27663 57443
rect 27663 57409 27672 57443
rect 27620 57400 27672 57409
rect 30012 57400 30064 57452
rect 33876 57477 33885 57511
rect 33885 57477 33919 57511
rect 33919 57477 33928 57511
rect 33876 57468 33928 57477
rect 37648 57511 37700 57520
rect 37648 57477 37657 57511
rect 37657 57477 37691 57511
rect 37691 57477 37700 57511
rect 37648 57468 37700 57477
rect 38752 57468 38804 57520
rect 24216 57332 24268 57384
rect 28080 57332 28132 57384
rect 30380 57332 30432 57384
rect 31576 57332 31628 57384
rect 32588 57443 32640 57452
rect 32588 57409 32597 57443
rect 32597 57409 32631 57443
rect 32631 57409 32640 57443
rect 32588 57400 32640 57409
rect 32864 57400 32916 57452
rect 33692 57443 33744 57452
rect 15752 57264 15804 57273
rect 26240 57307 26292 57316
rect 17960 57196 18012 57248
rect 26240 57273 26249 57307
rect 26249 57273 26283 57307
rect 26283 57273 26292 57307
rect 26240 57264 26292 57273
rect 31300 57264 31352 57316
rect 33692 57409 33701 57443
rect 33701 57409 33735 57443
rect 33735 57409 33744 57443
rect 33692 57400 33744 57409
rect 36084 57443 36136 57452
rect 36084 57409 36093 57443
rect 36093 57409 36127 57443
rect 36127 57409 36136 57443
rect 36084 57400 36136 57409
rect 37372 57400 37424 57452
rect 38844 57443 38896 57452
rect 34520 57375 34572 57384
rect 34520 57341 34529 57375
rect 34529 57341 34563 57375
rect 34563 57341 34572 57375
rect 34520 57332 34572 57341
rect 37648 57332 37700 57384
rect 38844 57409 38853 57443
rect 38853 57409 38887 57443
rect 38887 57409 38896 57443
rect 38844 57400 38896 57409
rect 41328 57443 41380 57452
rect 41328 57409 41337 57443
rect 41337 57409 41371 57443
rect 41371 57409 41380 57443
rect 41328 57400 41380 57409
rect 42984 57400 43036 57452
rect 43720 57400 43772 57452
rect 46388 57400 46440 57452
rect 53104 57400 53156 57452
rect 66996 57400 67048 57452
rect 38660 57332 38712 57384
rect 39120 57332 39172 57384
rect 42800 57375 42852 57384
rect 42800 57341 42809 57375
rect 42809 57341 42843 57375
rect 42843 57341 42852 57375
rect 42800 57332 42852 57341
rect 42892 57375 42944 57384
rect 42892 57341 42901 57375
rect 42901 57341 42935 57375
rect 42935 57341 42944 57375
rect 42892 57332 42944 57341
rect 35900 57264 35952 57316
rect 36176 57264 36228 57316
rect 19248 57196 19300 57248
rect 22376 57196 22428 57248
rect 30196 57196 30248 57248
rect 34152 57196 34204 57248
rect 38936 57196 38988 57248
rect 41144 57239 41196 57248
rect 41144 57205 41153 57239
rect 41153 57205 41187 57239
rect 41187 57205 41196 57239
rect 41144 57196 41196 57205
rect 42616 57196 42668 57248
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 65654 57094 65706 57146
rect 65718 57094 65770 57146
rect 65782 57094 65834 57146
rect 65846 57094 65898 57146
rect 65910 57094 65962 57146
rect 14372 57035 14424 57044
rect 14372 57001 14381 57035
rect 14381 57001 14415 57035
rect 14415 57001 14424 57035
rect 14372 56992 14424 57001
rect 23204 56992 23256 57044
rect 24216 56992 24268 57044
rect 28724 56992 28776 57044
rect 33968 57035 34020 57044
rect 33968 57001 33977 57035
rect 33977 57001 34011 57035
rect 34011 57001 34020 57035
rect 33968 56992 34020 57001
rect 37648 57035 37700 57044
rect 37648 57001 37657 57035
rect 37657 57001 37691 57035
rect 37691 57001 37700 57035
rect 37648 56992 37700 57001
rect 38844 56992 38896 57044
rect 42892 56992 42944 57044
rect 30380 56924 30432 56976
rect 34796 56924 34848 56976
rect 35348 56967 35400 56976
rect 35348 56933 35357 56967
rect 35357 56933 35391 56967
rect 35391 56933 35400 56967
rect 35348 56924 35400 56933
rect 15752 56856 15804 56908
rect 1400 56831 1452 56840
rect 1400 56797 1409 56831
rect 1409 56797 1443 56831
rect 1443 56797 1452 56831
rect 1400 56788 1452 56797
rect 13820 56788 13872 56840
rect 15200 56831 15252 56840
rect 15200 56797 15209 56831
rect 15209 56797 15243 56831
rect 15243 56797 15252 56831
rect 15200 56788 15252 56797
rect 36268 56899 36320 56908
rect 36268 56865 36277 56899
rect 36277 56865 36311 56899
rect 36311 56865 36320 56899
rect 36268 56856 36320 56865
rect 40776 56899 40828 56908
rect 40776 56865 40785 56899
rect 40785 56865 40819 56899
rect 40819 56865 40828 56899
rect 40776 56856 40828 56865
rect 43076 56899 43128 56908
rect 43076 56865 43085 56899
rect 43085 56865 43119 56899
rect 43119 56865 43128 56899
rect 43076 56856 43128 56865
rect 18144 56831 18196 56840
rect 18144 56797 18153 56831
rect 18153 56797 18187 56831
rect 18187 56797 18196 56831
rect 18144 56788 18196 56797
rect 18236 56831 18288 56840
rect 18236 56797 18245 56831
rect 18245 56797 18279 56831
rect 18279 56797 18288 56831
rect 18236 56788 18288 56797
rect 19432 56788 19484 56840
rect 19984 56788 20036 56840
rect 20536 56831 20588 56840
rect 20536 56797 20545 56831
rect 20545 56797 20579 56831
rect 20579 56797 20588 56831
rect 20536 56788 20588 56797
rect 21732 56788 21784 56840
rect 22192 56788 22244 56840
rect 26148 56831 26200 56840
rect 26148 56797 26157 56831
rect 26157 56797 26191 56831
rect 26191 56797 26200 56831
rect 26148 56788 26200 56797
rect 30840 56831 30892 56840
rect 30840 56797 30849 56831
rect 30849 56797 30883 56831
rect 30883 56797 30892 56831
rect 30840 56788 30892 56797
rect 34152 56831 34204 56840
rect 25044 56720 25096 56772
rect 26516 56720 26568 56772
rect 28632 56720 28684 56772
rect 31392 56720 31444 56772
rect 34152 56797 34161 56831
rect 34161 56797 34195 56831
rect 34195 56797 34204 56831
rect 34152 56788 34204 56797
rect 36544 56831 36596 56840
rect 36544 56797 36578 56831
rect 36578 56797 36596 56831
rect 36544 56788 36596 56797
rect 38936 56831 38988 56840
rect 38936 56797 38945 56831
rect 38945 56797 38979 56831
rect 38979 56797 38988 56831
rect 38936 56788 38988 56797
rect 42524 56788 42576 56840
rect 45376 56831 45428 56840
rect 45376 56797 45385 56831
rect 45385 56797 45419 56831
rect 45419 56797 45428 56831
rect 45376 56788 45428 56797
rect 46848 56831 46900 56840
rect 46848 56797 46857 56831
rect 46857 56797 46891 56831
rect 46891 56797 46900 56831
rect 46848 56788 46900 56797
rect 50620 56788 50672 56840
rect 67548 56788 67600 56840
rect 35072 56720 35124 56772
rect 35348 56720 35400 56772
rect 38200 56720 38252 56772
rect 41144 56720 41196 56772
rect 43352 56763 43404 56772
rect 43352 56729 43386 56763
rect 43386 56729 43404 56763
rect 43352 56720 43404 56729
rect 47584 56720 47636 56772
rect 1492 56652 1544 56704
rect 15384 56695 15436 56704
rect 15384 56661 15393 56695
rect 15393 56661 15427 56695
rect 15427 56661 15436 56695
rect 15384 56652 15436 56661
rect 16948 56695 17000 56704
rect 16948 56661 16957 56695
rect 16957 56661 16991 56695
rect 16991 56661 17000 56695
rect 16948 56652 17000 56661
rect 19432 56652 19484 56704
rect 20352 56695 20404 56704
rect 20352 56661 20361 56695
rect 20361 56661 20395 56695
rect 20395 56661 20404 56695
rect 20352 56652 20404 56661
rect 22192 56652 22244 56704
rect 27528 56695 27580 56704
rect 27528 56661 27537 56695
rect 27537 56661 27571 56695
rect 27571 56661 27580 56695
rect 27528 56652 27580 56661
rect 30380 56652 30432 56704
rect 33324 56695 33376 56704
rect 33324 56661 33333 56695
rect 33333 56661 33367 56695
rect 33367 56661 33376 56695
rect 33324 56652 33376 56661
rect 38752 56695 38804 56704
rect 38752 56661 38761 56695
rect 38761 56661 38795 56695
rect 38795 56661 38804 56695
rect 38752 56652 38804 56661
rect 38844 56695 38896 56704
rect 38844 56661 38853 56695
rect 38853 56661 38887 56695
rect 38887 56661 38896 56695
rect 38844 56652 38896 56661
rect 40500 56652 40552 56704
rect 42156 56695 42208 56704
rect 42156 56661 42165 56695
rect 42165 56661 42199 56695
rect 42199 56661 42208 56695
rect 42156 56652 42208 56661
rect 45192 56652 45244 56704
rect 48228 56695 48280 56704
rect 48228 56661 48237 56695
rect 48237 56661 48271 56695
rect 48271 56661 48280 56695
rect 48228 56652 48280 56661
rect 50160 56695 50212 56704
rect 50160 56661 50169 56695
rect 50169 56661 50203 56695
rect 50203 56661 50212 56695
rect 50160 56652 50212 56661
rect 67088 56652 67140 56704
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 2136 56448 2188 56500
rect 26148 56491 26200 56500
rect 16948 56423 17000 56432
rect 16948 56389 16982 56423
rect 16982 56389 17000 56423
rect 16948 56380 17000 56389
rect 20352 56380 20404 56432
rect 26148 56457 26157 56491
rect 26157 56457 26191 56491
rect 26191 56457 26200 56491
rect 26148 56448 26200 56457
rect 28540 56448 28592 56500
rect 29644 56448 29696 56500
rect 30932 56448 30984 56500
rect 35072 56448 35124 56500
rect 37372 56448 37424 56500
rect 40684 56448 40736 56500
rect 41328 56448 41380 56500
rect 43352 56491 43404 56500
rect 43352 56457 43361 56491
rect 43361 56457 43395 56491
rect 43395 56457 43404 56491
rect 43352 56448 43404 56457
rect 26884 56380 26936 56432
rect 27528 56380 27580 56432
rect 15384 56312 15436 56364
rect 19432 56312 19484 56364
rect 21732 56312 21784 56364
rect 22192 56355 22244 56364
rect 22192 56321 22201 56355
rect 22201 56321 22235 56355
rect 22235 56321 22244 56355
rect 22192 56312 22244 56321
rect 22376 56312 22428 56364
rect 24952 56312 25004 56364
rect 25412 56312 25464 56364
rect 26424 56312 26476 56364
rect 28540 56312 28592 56364
rect 33324 56380 33376 56432
rect 36728 56380 36780 56432
rect 16028 56244 16080 56296
rect 27160 56287 27212 56296
rect 27160 56253 27169 56287
rect 27169 56253 27203 56287
rect 27203 56253 27212 56287
rect 27160 56244 27212 56253
rect 14924 56219 14976 56228
rect 14924 56185 14933 56219
rect 14933 56185 14967 56219
rect 14967 56185 14976 56219
rect 14924 56176 14976 56185
rect 18144 56176 18196 56228
rect 28448 56176 28500 56228
rect 19340 56108 19392 56160
rect 22744 56108 22796 56160
rect 24492 56108 24544 56160
rect 25320 56151 25372 56160
rect 25320 56117 25329 56151
rect 25329 56117 25363 56151
rect 25363 56117 25372 56151
rect 25320 56108 25372 56117
rect 30104 56244 30156 56296
rect 30196 56287 30248 56296
rect 30196 56253 30205 56287
rect 30205 56253 30239 56287
rect 30239 56253 30248 56287
rect 30196 56244 30248 56253
rect 33048 56244 33100 56296
rect 36176 56312 36228 56364
rect 37372 56312 37424 56364
rect 38752 56312 38804 56364
rect 40500 56355 40552 56364
rect 35992 56244 36044 56296
rect 37188 56244 37240 56296
rect 38844 56244 38896 56296
rect 40500 56321 40509 56355
rect 40509 56321 40543 56355
rect 40543 56321 40552 56355
rect 40500 56312 40552 56321
rect 40684 56355 40736 56364
rect 40684 56321 40693 56355
rect 40693 56321 40727 56355
rect 40727 56321 40736 56355
rect 40684 56312 40736 56321
rect 42892 56380 42944 56432
rect 50160 56380 50212 56432
rect 43536 56355 43588 56364
rect 43536 56321 43545 56355
rect 43545 56321 43579 56355
rect 43579 56321 43588 56355
rect 43536 56312 43588 56321
rect 45192 56355 45244 56364
rect 45192 56321 45201 56355
rect 45201 56321 45235 56355
rect 45235 56321 45244 56355
rect 45192 56312 45244 56321
rect 45836 56312 45888 56364
rect 48228 56355 48280 56364
rect 48228 56321 48237 56355
rect 48237 56321 48271 56355
rect 48271 56321 48280 56355
rect 48228 56312 48280 56321
rect 49700 56312 49752 56364
rect 50344 56312 50396 56364
rect 29644 56219 29696 56228
rect 29644 56185 29653 56219
rect 29653 56185 29687 56219
rect 29687 56185 29696 56219
rect 29644 56176 29696 56185
rect 34612 56176 34664 56228
rect 36636 56176 36688 56228
rect 38200 56176 38252 56228
rect 41604 56176 41656 56228
rect 42156 56244 42208 56296
rect 42800 56244 42852 56296
rect 43904 56244 43956 56296
rect 48780 56244 48832 56296
rect 42616 56176 42668 56228
rect 30380 56108 30432 56160
rect 32312 56108 32364 56160
rect 35808 56108 35860 56160
rect 35900 56108 35952 56160
rect 37096 56108 37148 56160
rect 42432 56151 42484 56160
rect 42432 56117 42441 56151
rect 42441 56117 42475 56151
rect 42475 56117 42484 56151
rect 42432 56108 42484 56117
rect 42984 56108 43036 56160
rect 46572 56151 46624 56160
rect 46572 56117 46581 56151
rect 46581 56117 46615 56151
rect 46615 56117 46624 56151
rect 46572 56108 46624 56117
rect 47768 56108 47820 56160
rect 50528 56151 50580 56160
rect 50528 56117 50537 56151
rect 50537 56117 50571 56151
rect 50571 56117 50580 56151
rect 50528 56108 50580 56117
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 65654 56006 65706 56058
rect 65718 56006 65770 56058
rect 65782 56006 65834 56058
rect 65846 56006 65898 56058
rect 65910 56006 65962 56058
rect 16028 55947 16080 55956
rect 16028 55913 16037 55947
rect 16037 55913 16071 55947
rect 16071 55913 16080 55947
rect 16028 55904 16080 55913
rect 20536 55904 20588 55956
rect 22836 55904 22888 55956
rect 26516 55947 26568 55956
rect 26516 55913 26525 55947
rect 26525 55913 26559 55947
rect 26559 55913 26568 55947
rect 26516 55904 26568 55913
rect 26884 55904 26936 55956
rect 20444 55836 20496 55888
rect 30012 55836 30064 55888
rect 30288 55904 30340 55956
rect 30840 55904 30892 55956
rect 34612 55836 34664 55888
rect 24492 55811 24544 55820
rect 24492 55777 24501 55811
rect 24501 55777 24535 55811
rect 24535 55777 24544 55811
rect 24492 55768 24544 55777
rect 15292 55700 15344 55752
rect 17316 55700 17368 55752
rect 23204 55700 23256 55752
rect 25320 55700 25372 55752
rect 28448 55811 28500 55820
rect 28448 55777 28457 55811
rect 28457 55777 28491 55811
rect 28491 55777 28500 55811
rect 28448 55768 28500 55777
rect 19340 55632 19392 55684
rect 22192 55632 22244 55684
rect 27620 55700 27672 55752
rect 28356 55700 28408 55752
rect 34796 55768 34848 55820
rect 29828 55700 29880 55752
rect 30564 55700 30616 55752
rect 32312 55743 32364 55752
rect 32312 55709 32321 55743
rect 32321 55709 32355 55743
rect 32355 55709 32364 55743
rect 32312 55700 32364 55709
rect 36820 55904 36872 55956
rect 45836 55947 45888 55956
rect 45836 55913 45845 55947
rect 45845 55913 45879 55947
rect 45879 55913 45888 55947
rect 45836 55904 45888 55913
rect 46848 55947 46900 55956
rect 46848 55913 46857 55947
rect 46857 55913 46891 55947
rect 46891 55913 46900 55947
rect 46848 55904 46900 55913
rect 46940 55904 46992 55956
rect 48596 55904 48648 55956
rect 48780 55947 48832 55956
rect 48780 55913 48789 55947
rect 48789 55913 48823 55947
rect 48823 55913 48832 55947
rect 48780 55904 48832 55913
rect 50620 55904 50672 55956
rect 36084 55768 36136 55820
rect 36636 55768 36688 55820
rect 27528 55632 27580 55684
rect 14648 55607 14700 55616
rect 14648 55573 14657 55607
rect 14657 55573 14691 55607
rect 14691 55573 14700 55607
rect 14648 55564 14700 55573
rect 16948 55564 17000 55616
rect 20076 55607 20128 55616
rect 20076 55573 20101 55607
rect 20101 55573 20128 55607
rect 20076 55564 20128 55573
rect 25136 55564 25188 55616
rect 30104 55632 30156 55684
rect 30380 55675 30432 55684
rect 30380 55641 30389 55675
rect 30389 55641 30423 55675
rect 30423 55641 30432 55675
rect 30380 55632 30432 55641
rect 32680 55632 32732 55684
rect 34152 55675 34204 55684
rect 34152 55641 34161 55675
rect 34161 55641 34195 55675
rect 34195 55641 34204 55675
rect 34152 55632 34204 55641
rect 28724 55564 28776 55616
rect 29736 55564 29788 55616
rect 30472 55564 30524 55616
rect 30748 55607 30800 55616
rect 30748 55573 30757 55607
rect 30757 55573 30791 55607
rect 30791 55573 30800 55607
rect 30748 55564 30800 55573
rect 34612 55564 34664 55616
rect 36268 55700 36320 55752
rect 36820 55700 36872 55752
rect 37188 55700 37240 55752
rect 35900 55632 35952 55684
rect 38200 55743 38252 55752
rect 38200 55709 38209 55743
rect 38209 55709 38243 55743
rect 38243 55709 38252 55743
rect 38200 55700 38252 55709
rect 38752 55768 38804 55820
rect 39120 55768 39172 55820
rect 46572 55768 46624 55820
rect 55680 55836 55732 55888
rect 48228 55768 48280 55820
rect 38936 55743 38988 55752
rect 38936 55709 38945 55743
rect 38945 55709 38979 55743
rect 38979 55709 38988 55743
rect 38936 55700 38988 55709
rect 39028 55743 39080 55752
rect 39028 55709 39037 55743
rect 39037 55709 39071 55743
rect 39071 55709 39080 55743
rect 39028 55700 39080 55709
rect 36636 55564 36688 55616
rect 37188 55607 37240 55616
rect 37188 55573 37197 55607
rect 37197 55573 37231 55607
rect 37231 55573 37240 55607
rect 37188 55564 37240 55573
rect 38660 55607 38712 55616
rect 38660 55573 38669 55607
rect 38669 55573 38703 55607
rect 38703 55573 38712 55607
rect 38660 55564 38712 55573
rect 40776 55700 40828 55752
rect 45192 55743 45244 55752
rect 45192 55709 45201 55743
rect 45201 55709 45235 55743
rect 45235 55709 45244 55743
rect 45192 55700 45244 55709
rect 40500 55632 40552 55684
rect 46940 55700 46992 55752
rect 50528 55768 50580 55820
rect 48596 55743 48648 55752
rect 48596 55709 48605 55743
rect 48605 55709 48639 55743
rect 48639 55709 48648 55743
rect 50344 55743 50396 55752
rect 48596 55700 48648 55709
rect 50344 55709 50353 55743
rect 50353 55709 50387 55743
rect 50387 55709 50396 55743
rect 50344 55700 50396 55709
rect 47952 55564 48004 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 25412 55403 25464 55412
rect 25412 55369 25421 55403
rect 25421 55369 25455 55403
rect 25455 55369 25464 55403
rect 25412 55360 25464 55369
rect 27160 55360 27212 55412
rect 28540 55403 28592 55412
rect 28540 55369 28549 55403
rect 28549 55369 28583 55403
rect 28583 55369 28592 55403
rect 28540 55360 28592 55369
rect 31392 55403 31444 55412
rect 31392 55369 31401 55403
rect 31401 55369 31435 55403
rect 31435 55369 31444 55403
rect 31392 55360 31444 55369
rect 32680 55403 32732 55412
rect 32680 55369 32689 55403
rect 32689 55369 32723 55403
rect 32723 55369 32732 55403
rect 32680 55360 32732 55369
rect 36636 55403 36688 55412
rect 36636 55369 36645 55403
rect 36645 55369 36679 55403
rect 36679 55369 36688 55403
rect 36636 55360 36688 55369
rect 39028 55360 39080 55412
rect 40500 55403 40552 55412
rect 40500 55369 40509 55403
rect 40509 55369 40543 55403
rect 40543 55369 40552 55403
rect 40500 55360 40552 55369
rect 43904 55403 43956 55412
rect 43904 55369 43913 55403
rect 43913 55369 43947 55403
rect 43947 55369 43956 55403
rect 43904 55360 43956 55369
rect 47584 55403 47636 55412
rect 47584 55369 47593 55403
rect 47593 55369 47627 55403
rect 47627 55369 47636 55403
rect 47584 55360 47636 55369
rect 14648 55292 14700 55344
rect 13820 55224 13872 55276
rect 16948 55267 17000 55276
rect 16948 55233 16957 55267
rect 16957 55233 16991 55267
rect 16991 55233 17000 55267
rect 16948 55224 17000 55233
rect 17684 55224 17736 55276
rect 18236 55224 18288 55276
rect 22928 55224 22980 55276
rect 25136 55267 25188 55276
rect 25136 55233 25145 55267
rect 25145 55233 25179 55267
rect 25179 55233 25188 55267
rect 25136 55224 25188 55233
rect 25504 55224 25556 55276
rect 15568 55063 15620 55072
rect 15568 55029 15577 55063
rect 15577 55029 15611 55063
rect 15611 55029 15620 55063
rect 15568 55020 15620 55029
rect 18052 55020 18104 55072
rect 25688 55224 25740 55276
rect 28724 55267 28776 55276
rect 28724 55233 28733 55267
rect 28733 55233 28767 55267
rect 28767 55233 28776 55267
rect 28724 55224 28776 55233
rect 30748 55224 30800 55276
rect 32220 55224 32272 55276
rect 32496 55224 32548 55276
rect 33048 55224 33100 55276
rect 34704 55224 34756 55276
rect 35532 55224 35584 55276
rect 36268 55292 36320 55344
rect 36728 55292 36780 55344
rect 36084 55224 36136 55276
rect 37188 55224 37240 55276
rect 39120 55267 39172 55276
rect 39120 55233 39129 55267
rect 39129 55233 39163 55267
rect 39163 55233 39172 55267
rect 39120 55224 39172 55233
rect 41328 55224 41380 55276
rect 42524 55267 42576 55276
rect 42524 55233 42533 55267
rect 42533 55233 42567 55267
rect 42567 55233 42576 55267
rect 42524 55224 42576 55233
rect 43168 55224 43220 55276
rect 45836 55267 45888 55276
rect 45836 55233 45845 55267
rect 45845 55233 45879 55267
rect 45879 55233 45888 55267
rect 45836 55224 45888 55233
rect 47768 55267 47820 55276
rect 47768 55233 47777 55267
rect 47777 55233 47811 55267
rect 47811 55233 47820 55267
rect 47768 55224 47820 55233
rect 48504 55267 48556 55276
rect 48504 55233 48513 55267
rect 48513 55233 48547 55267
rect 48547 55233 48556 55267
rect 48504 55224 48556 55233
rect 51264 55267 51316 55276
rect 51264 55233 51273 55267
rect 51273 55233 51307 55267
rect 51307 55233 51316 55267
rect 51264 55224 51316 55233
rect 39028 55156 39080 55208
rect 42432 55156 42484 55208
rect 35992 55088 36044 55140
rect 36268 55088 36320 55140
rect 19156 55063 19208 55072
rect 19156 55029 19165 55063
rect 19165 55029 19199 55063
rect 19199 55029 19208 55063
rect 19156 55020 19208 55029
rect 35440 55020 35492 55072
rect 35808 55063 35860 55072
rect 35808 55029 35817 55063
rect 35817 55029 35851 55063
rect 35851 55029 35860 55063
rect 35808 55020 35860 55029
rect 37832 55063 37884 55072
rect 37832 55029 37841 55063
rect 37841 55029 37875 55063
rect 37875 55029 37884 55063
rect 37832 55020 37884 55029
rect 45744 55063 45796 55072
rect 45744 55029 45753 55063
rect 45753 55029 45787 55063
rect 45787 55029 45796 55063
rect 45744 55020 45796 55029
rect 48320 55063 48372 55072
rect 48320 55029 48329 55063
rect 48329 55029 48363 55063
rect 48363 55029 48372 55063
rect 48320 55020 48372 55029
rect 50436 55020 50488 55072
rect 51080 55063 51132 55072
rect 51080 55029 51089 55063
rect 51089 55029 51123 55063
rect 51123 55029 51132 55063
rect 51080 55020 51132 55029
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 65654 54918 65706 54970
rect 65718 54918 65770 54970
rect 65782 54918 65834 54970
rect 65846 54918 65898 54970
rect 65910 54918 65962 54970
rect 15292 54859 15344 54868
rect 15292 54825 15301 54859
rect 15301 54825 15335 54859
rect 15335 54825 15344 54859
rect 15292 54816 15344 54825
rect 17684 54859 17736 54868
rect 17684 54825 17693 54859
rect 17693 54825 17727 54859
rect 17727 54825 17736 54859
rect 17684 54816 17736 54825
rect 22192 54816 22244 54868
rect 34704 54859 34756 54868
rect 34704 54825 34713 54859
rect 34713 54825 34747 54859
rect 34747 54825 34756 54859
rect 34704 54816 34756 54825
rect 35716 54816 35768 54868
rect 38660 54859 38712 54868
rect 21824 54748 21876 54800
rect 15200 54612 15252 54664
rect 19156 54612 19208 54664
rect 19984 54612 20036 54664
rect 20352 54655 20404 54664
rect 20352 54621 20361 54655
rect 20361 54621 20395 54655
rect 20395 54621 20404 54655
rect 20352 54612 20404 54621
rect 21732 54680 21784 54732
rect 22836 54748 22888 54800
rect 33324 54748 33376 54800
rect 15568 54544 15620 54596
rect 18236 54544 18288 54596
rect 19248 54544 19300 54596
rect 17500 54476 17552 54528
rect 19340 54476 19392 54528
rect 19432 54476 19484 54528
rect 20168 54519 20220 54528
rect 20168 54485 20177 54519
rect 20177 54485 20211 54519
rect 20211 54485 20220 54519
rect 20168 54476 20220 54485
rect 21916 54544 21968 54596
rect 22836 54612 22888 54664
rect 24032 54680 24084 54732
rect 23388 54655 23440 54664
rect 23388 54621 23397 54655
rect 23397 54621 23431 54655
rect 23431 54621 23440 54655
rect 23388 54612 23440 54621
rect 25412 54655 25464 54664
rect 23020 54544 23072 54596
rect 25412 54621 25421 54655
rect 25421 54621 25455 54655
rect 25455 54621 25464 54655
rect 25412 54612 25464 54621
rect 29000 54655 29052 54664
rect 29000 54621 29009 54655
rect 29009 54621 29043 54655
rect 29043 54621 29052 54655
rect 29000 54612 29052 54621
rect 30564 54612 30616 54664
rect 31668 54680 31720 54732
rect 31760 54655 31812 54664
rect 31760 54621 31769 54655
rect 31769 54621 31803 54655
rect 31803 54621 31812 54655
rect 31760 54612 31812 54621
rect 31852 54655 31904 54664
rect 31852 54621 31861 54655
rect 31861 54621 31895 54655
rect 31895 54621 31904 54655
rect 31852 54612 31904 54621
rect 35440 54612 35492 54664
rect 35716 54612 35768 54664
rect 38660 54825 38669 54859
rect 38669 54825 38703 54859
rect 38703 54825 38712 54859
rect 38660 54816 38712 54825
rect 41328 54680 41380 54732
rect 45376 54816 45428 54868
rect 46940 54816 46992 54868
rect 45744 54723 45796 54732
rect 38936 54612 38988 54664
rect 43076 54612 43128 54664
rect 45744 54689 45753 54723
rect 45753 54689 45787 54723
rect 45787 54689 45796 54723
rect 45744 54680 45796 54689
rect 50436 54723 50488 54732
rect 50436 54689 50445 54723
rect 50445 54689 50479 54723
rect 50479 54689 50488 54723
rect 50436 54680 50488 54689
rect 45008 54655 45060 54664
rect 45008 54621 45017 54655
rect 45017 54621 45051 54655
rect 45051 54621 45060 54655
rect 45008 54612 45060 54621
rect 47676 54655 47728 54664
rect 47676 54621 47685 54655
rect 47685 54621 47719 54655
rect 47719 54621 47728 54655
rect 47676 54612 47728 54621
rect 48320 54612 48372 54664
rect 51080 54612 51132 54664
rect 30012 54544 30064 54596
rect 32404 54587 32456 54596
rect 32404 54553 32413 54587
rect 32413 54553 32447 54587
rect 32447 54553 32456 54587
rect 32404 54544 32456 54553
rect 22284 54476 22336 54528
rect 23296 54476 23348 54528
rect 25136 54476 25188 54528
rect 29828 54476 29880 54528
rect 36728 54544 36780 54596
rect 41420 54544 41472 54596
rect 41604 54544 41656 54596
rect 43168 54587 43220 54596
rect 43168 54553 43177 54587
rect 43177 54553 43211 54587
rect 43211 54553 43220 54587
rect 43168 54544 43220 54553
rect 45652 54544 45704 54596
rect 38108 54476 38160 54528
rect 38292 54519 38344 54528
rect 38292 54485 38301 54519
rect 38301 54485 38335 54519
rect 38335 54485 38344 54519
rect 38292 54476 38344 54485
rect 43628 54476 43680 54528
rect 46572 54476 46624 54528
rect 48688 54476 48740 54528
rect 49884 54476 49936 54528
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 33140 54272 33192 54324
rect 19248 54204 19300 54256
rect 20168 54204 20220 54256
rect 21916 54204 21968 54256
rect 22192 54247 22244 54256
rect 22192 54213 22201 54247
rect 22201 54213 22235 54247
rect 22235 54213 22244 54247
rect 22192 54204 22244 54213
rect 16580 54136 16632 54188
rect 6552 54111 6604 54120
rect 6552 54077 6561 54111
rect 6561 54077 6595 54111
rect 6595 54077 6604 54111
rect 6552 54068 6604 54077
rect 17500 54111 17552 54120
rect 3516 54000 3568 54052
rect 17500 54077 17509 54111
rect 17509 54077 17543 54111
rect 17543 54077 17552 54111
rect 17500 54068 17552 54077
rect 18236 54179 18288 54188
rect 18236 54145 18245 54179
rect 18245 54145 18279 54179
rect 18279 54145 18288 54179
rect 18236 54136 18288 54145
rect 19432 54136 19484 54188
rect 21732 54136 21784 54188
rect 29000 54204 29052 54256
rect 23204 54179 23256 54188
rect 18052 54068 18104 54120
rect 18328 54111 18380 54120
rect 18328 54077 18362 54111
rect 18362 54077 18380 54111
rect 18328 54068 18380 54077
rect 18512 54111 18564 54120
rect 18512 54077 18521 54111
rect 18521 54077 18555 54111
rect 18555 54077 18564 54111
rect 18512 54068 18564 54077
rect 20628 54068 20680 54120
rect 23204 54145 23213 54179
rect 23213 54145 23247 54179
rect 23247 54145 23256 54179
rect 23204 54136 23256 54145
rect 23296 54136 23348 54188
rect 24952 54136 25004 54188
rect 26332 54179 26384 54188
rect 26332 54145 26341 54179
rect 26341 54145 26375 54179
rect 26375 54145 26384 54179
rect 26332 54136 26384 54145
rect 27068 54136 27120 54188
rect 29828 54179 29880 54188
rect 29828 54145 29837 54179
rect 29837 54145 29871 54179
rect 29871 54145 29880 54179
rect 29828 54136 29880 54145
rect 30656 54136 30708 54188
rect 38292 54204 38344 54256
rect 45192 54272 45244 54324
rect 45652 54315 45704 54324
rect 45652 54281 45661 54315
rect 45661 54281 45695 54315
rect 45695 54281 45704 54315
rect 45652 54272 45704 54281
rect 47676 54272 47728 54324
rect 48504 54272 48556 54324
rect 51264 54272 51316 54324
rect 32864 54136 32916 54188
rect 37556 54179 37608 54188
rect 37556 54145 37565 54179
rect 37565 54145 37599 54179
rect 37599 54145 37608 54179
rect 37556 54136 37608 54145
rect 40040 54179 40092 54188
rect 40040 54145 40049 54179
rect 40049 54145 40083 54179
rect 40083 54145 40092 54179
rect 40040 54136 40092 54145
rect 41420 54179 41472 54188
rect 41420 54145 41429 54179
rect 41429 54145 41463 54179
rect 41463 54145 41472 54179
rect 41420 54136 41472 54145
rect 17960 54043 18012 54052
rect 17960 54009 17969 54043
rect 17969 54009 18003 54043
rect 18003 54009 18012 54043
rect 17960 54000 18012 54009
rect 1952 53975 2004 53984
rect 1952 53941 1961 53975
rect 1961 53941 1995 53975
rect 1995 53941 2004 53975
rect 1952 53932 2004 53941
rect 16856 53932 16908 53984
rect 16948 53932 17000 53984
rect 18328 53932 18380 53984
rect 19340 53932 19392 53984
rect 22836 53932 22888 53984
rect 24860 53932 24912 53984
rect 29184 54000 29236 54052
rect 28356 53975 28408 53984
rect 28356 53941 28365 53975
rect 28365 53941 28399 53975
rect 28399 53941 28408 53975
rect 28356 53932 28408 53941
rect 29828 53932 29880 53984
rect 32772 53932 32824 53984
rect 37832 53932 37884 53984
rect 41328 54000 41380 54052
rect 43628 54179 43680 54188
rect 43628 54145 43637 54179
rect 43637 54145 43671 54179
rect 43671 54145 43680 54179
rect 43628 54136 43680 54145
rect 43720 54136 43772 54188
rect 46940 54136 46992 54188
rect 48688 54179 48740 54188
rect 48688 54145 48697 54179
rect 48697 54145 48731 54179
rect 48731 54145 48740 54179
rect 48688 54136 48740 54145
rect 49700 54136 49752 54188
rect 50068 54179 50120 54188
rect 50068 54145 50077 54179
rect 50077 54145 50111 54179
rect 50111 54145 50120 54179
rect 50068 54136 50120 54145
rect 50160 54136 50212 54188
rect 46572 54068 46624 54120
rect 49884 54111 49936 54120
rect 49884 54077 49893 54111
rect 49893 54077 49927 54111
rect 49927 54077 49936 54111
rect 49884 54068 49936 54077
rect 38936 53975 38988 53984
rect 38936 53941 38945 53975
rect 38945 53941 38979 53975
rect 38979 53941 38988 53975
rect 38936 53932 38988 53941
rect 40776 53975 40828 53984
rect 40776 53941 40785 53975
rect 40785 53941 40819 53975
rect 40819 53941 40828 53975
rect 40776 53932 40828 53941
rect 41512 53975 41564 53984
rect 41512 53941 41521 53975
rect 41521 53941 41555 53975
rect 41555 53941 41564 53975
rect 41512 53932 41564 53941
rect 45468 53932 45520 53984
rect 45560 53932 45612 53984
rect 50804 53932 50856 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 65654 53830 65706 53882
rect 65718 53830 65770 53882
rect 65782 53830 65834 53882
rect 65846 53830 65898 53882
rect 65910 53830 65962 53882
rect 6552 53728 6604 53780
rect 16948 53771 17000 53780
rect 16948 53737 16957 53771
rect 16957 53737 16991 53771
rect 16991 53737 17000 53771
rect 16948 53728 17000 53737
rect 20352 53728 20404 53780
rect 23388 53728 23440 53780
rect 27068 53728 27120 53780
rect 27252 53728 27304 53780
rect 30012 53771 30064 53780
rect 20444 53660 20496 53712
rect 26240 53703 26292 53712
rect 26240 53669 26249 53703
rect 26249 53669 26283 53703
rect 26283 53669 26292 53703
rect 26240 53660 26292 53669
rect 29092 53660 29144 53712
rect 1952 53592 2004 53644
rect 2780 53635 2832 53644
rect 2780 53601 2789 53635
rect 2789 53601 2823 53635
rect 2823 53601 2832 53635
rect 2780 53592 2832 53601
rect 6368 53524 6420 53576
rect 13820 53524 13872 53576
rect 15200 53592 15252 53644
rect 22192 53592 22244 53644
rect 24860 53635 24912 53644
rect 24860 53601 24869 53635
rect 24869 53601 24903 53635
rect 24903 53601 24912 53635
rect 24860 53592 24912 53601
rect 15568 53567 15620 53576
rect 2412 53456 2464 53508
rect 15568 53533 15577 53567
rect 15577 53533 15611 53567
rect 15611 53533 15620 53567
rect 15568 53524 15620 53533
rect 17408 53567 17460 53576
rect 17408 53533 17417 53567
rect 17417 53533 17451 53567
rect 17451 53533 17460 53567
rect 17408 53524 17460 53533
rect 21732 53567 21784 53576
rect 15200 53456 15252 53508
rect 16672 53456 16724 53508
rect 18880 53456 18932 53508
rect 19340 53456 19392 53508
rect 21732 53533 21741 53567
rect 21741 53533 21775 53567
rect 21775 53533 21784 53567
rect 21732 53524 21784 53533
rect 20076 53456 20128 53508
rect 20168 53456 20220 53508
rect 25136 53567 25188 53576
rect 25136 53533 25170 53567
rect 25170 53533 25188 53567
rect 22192 53456 22244 53508
rect 13544 53388 13596 53440
rect 14280 53388 14332 53440
rect 17316 53388 17368 53440
rect 18604 53431 18656 53440
rect 18604 53397 18613 53431
rect 18613 53397 18647 53431
rect 18647 53397 18656 53431
rect 18604 53388 18656 53397
rect 25136 53524 25188 53533
rect 30012 53737 30021 53771
rect 30021 53737 30055 53771
rect 30055 53737 30064 53771
rect 30012 53728 30064 53737
rect 30288 53728 30340 53780
rect 30656 53771 30708 53780
rect 30656 53737 30665 53771
rect 30665 53737 30699 53771
rect 30699 53737 30708 53771
rect 30656 53728 30708 53737
rect 32864 53771 32916 53780
rect 32864 53737 32873 53771
rect 32873 53737 32907 53771
rect 32907 53737 32916 53771
rect 32864 53728 32916 53737
rect 37464 53728 37516 53780
rect 43536 53728 43588 53780
rect 43720 53728 43772 53780
rect 45836 53728 45888 53780
rect 47584 53728 47636 53780
rect 48688 53771 48740 53780
rect 48688 53737 48697 53771
rect 48697 53737 48731 53771
rect 48731 53737 48740 53771
rect 48688 53728 48740 53737
rect 30104 53660 30156 53712
rect 22560 53456 22612 53508
rect 27252 53456 27304 53508
rect 27804 53567 27856 53576
rect 27804 53533 27813 53567
rect 27813 53533 27847 53567
rect 27847 53533 27856 53567
rect 27804 53524 27856 53533
rect 29736 53524 29788 53576
rect 28356 53456 28408 53508
rect 29828 53499 29880 53508
rect 29828 53465 29837 53499
rect 29837 53465 29871 53499
rect 29871 53465 29880 53499
rect 29828 53456 29880 53465
rect 31760 53592 31812 53644
rect 35440 53592 35492 53644
rect 30104 53388 30156 53440
rect 32404 53524 32456 53576
rect 33140 53567 33192 53576
rect 33140 53533 33149 53567
rect 33149 53533 33183 53567
rect 33183 53533 33192 53567
rect 33140 53524 33192 53533
rect 33324 53567 33376 53576
rect 33324 53533 33333 53567
rect 33333 53533 33367 53567
rect 33367 53533 33376 53567
rect 33324 53524 33376 53533
rect 35256 53567 35308 53576
rect 34428 53456 34480 53508
rect 35256 53533 35265 53567
rect 35265 53533 35299 53567
rect 35299 53533 35308 53567
rect 35256 53524 35308 53533
rect 35624 53524 35676 53576
rect 35992 53524 36044 53576
rect 35716 53456 35768 53508
rect 35900 53388 35952 53440
rect 49884 53660 49936 53712
rect 41512 53635 41564 53644
rect 41512 53601 41521 53635
rect 41521 53601 41555 53635
rect 41555 53601 41564 53635
rect 41512 53592 41564 53601
rect 43168 53592 43220 53644
rect 37556 53524 37608 53576
rect 39396 53524 39448 53576
rect 41420 53524 41472 53576
rect 43720 53524 43772 53576
rect 45192 53592 45244 53644
rect 46572 53592 46624 53644
rect 37280 53456 37332 53508
rect 38844 53456 38896 53508
rect 40224 53456 40276 53508
rect 37924 53431 37976 53440
rect 37924 53397 37933 53431
rect 37933 53397 37967 53431
rect 37967 53397 37976 53431
rect 37924 53388 37976 53397
rect 39488 53388 39540 53440
rect 41788 53499 41840 53508
rect 41788 53465 41822 53499
rect 41822 53465 41840 53499
rect 41788 53456 41840 53465
rect 45008 53456 45060 53508
rect 46112 53524 46164 53576
rect 48504 53567 48556 53576
rect 48504 53533 48513 53567
rect 48513 53533 48547 53567
rect 48547 53533 48556 53567
rect 48504 53524 48556 53533
rect 50620 53524 50672 53576
rect 50804 53567 50856 53576
rect 50804 53533 50838 53567
rect 50838 53533 50856 53567
rect 50804 53524 50856 53533
rect 48228 53456 48280 53508
rect 42892 53431 42944 53440
rect 42892 53397 42901 53431
rect 42901 53397 42935 53431
rect 42935 53397 42944 53431
rect 42892 53388 42944 53397
rect 46204 53388 46256 53440
rect 46388 53431 46440 53440
rect 46388 53397 46397 53431
rect 46397 53397 46431 53431
rect 46431 53397 46440 53431
rect 46388 53388 46440 53397
rect 48964 53388 49016 53440
rect 49884 53388 49936 53440
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 2412 53227 2464 53236
rect 2412 53193 2421 53227
rect 2421 53193 2455 53227
rect 2455 53193 2464 53227
rect 2412 53184 2464 53193
rect 15568 53184 15620 53236
rect 16672 53227 16724 53236
rect 16672 53193 16681 53227
rect 16681 53193 16715 53227
rect 16715 53193 16724 53227
rect 16672 53184 16724 53193
rect 17408 53184 17460 53236
rect 22928 53184 22980 53236
rect 23296 53184 23348 53236
rect 25412 53184 25464 53236
rect 16764 53116 16816 53168
rect 24860 53116 24912 53168
rect 5172 53048 5224 53100
rect 13544 53091 13596 53100
rect 13544 53057 13553 53091
rect 13553 53057 13587 53091
rect 13587 53057 13596 53091
rect 13544 53048 13596 53057
rect 14096 53048 14148 53100
rect 15844 53048 15896 53100
rect 16856 53091 16908 53100
rect 16856 53057 16865 53091
rect 16865 53057 16899 53091
rect 16899 53057 16908 53091
rect 16856 53048 16908 53057
rect 19984 53048 20036 53100
rect 20904 53048 20956 53100
rect 21732 53048 21784 53100
rect 24400 53091 24452 53100
rect 24400 53057 24409 53091
rect 24409 53057 24443 53091
rect 24443 53057 24452 53091
rect 24400 53048 24452 53057
rect 26240 53116 26292 53168
rect 25504 53091 25556 53100
rect 25504 53057 25513 53091
rect 25513 53057 25547 53091
rect 25547 53057 25556 53091
rect 25504 53048 25556 53057
rect 22376 53023 22428 53032
rect 22376 52989 22385 53023
rect 22385 52989 22419 53023
rect 22419 52989 22428 53023
rect 22376 52980 22428 52989
rect 22560 52980 22612 53032
rect 26332 52980 26384 53032
rect 21732 52912 21784 52964
rect 24032 52912 24084 52964
rect 24492 52912 24544 52964
rect 31852 53184 31904 53236
rect 34796 53184 34848 53236
rect 35256 53184 35308 53236
rect 35900 53184 35952 53236
rect 37096 53184 37148 53236
rect 37280 53227 37332 53236
rect 37280 53193 37289 53227
rect 37289 53193 37323 53227
rect 37323 53193 37332 53227
rect 37280 53184 37332 53193
rect 40040 53184 40092 53236
rect 41236 53184 41288 53236
rect 41788 53227 41840 53236
rect 28448 53048 28500 53100
rect 29092 53091 29144 53100
rect 29092 53057 29126 53091
rect 29126 53057 29144 53091
rect 29092 53048 29144 53057
rect 28172 52980 28224 53032
rect 28356 52980 28408 53032
rect 29920 52980 29972 53032
rect 30748 52980 30800 53032
rect 35532 53116 35584 53168
rect 32496 53048 32548 53100
rect 33416 53091 33468 53100
rect 33416 53057 33450 53091
rect 33450 53057 33468 53091
rect 33416 53048 33468 53057
rect 35716 53048 35768 53100
rect 37464 53091 37516 53100
rect 1400 52844 1452 52896
rect 15200 52844 15252 52896
rect 16304 52844 16356 52896
rect 19340 52887 19392 52896
rect 19340 52853 19349 52887
rect 19349 52853 19383 52887
rect 19383 52853 19392 52887
rect 19340 52844 19392 52853
rect 22744 52844 22796 52896
rect 24584 52844 24636 52896
rect 27436 52887 27488 52896
rect 27436 52853 27445 52887
rect 27445 52853 27479 52887
rect 27479 52853 27488 52887
rect 27436 52844 27488 52853
rect 28816 52912 28868 52964
rect 29828 52844 29880 52896
rect 31208 52844 31260 52896
rect 32772 52980 32824 53032
rect 36084 53023 36136 53032
rect 31392 52912 31444 52964
rect 32680 52912 32732 52964
rect 36084 52989 36093 53023
rect 36093 52989 36127 53023
rect 36127 52989 36136 53023
rect 36084 52980 36136 52989
rect 37464 53057 37473 53091
rect 37473 53057 37507 53091
rect 37507 53057 37516 53091
rect 37464 53048 37516 53057
rect 37924 53116 37976 53168
rect 40776 53116 40828 53168
rect 41788 53193 41797 53227
rect 41797 53193 41831 53227
rect 41831 53193 41840 53227
rect 41788 53184 41840 53193
rect 42800 53184 42852 53236
rect 45560 53227 45612 53236
rect 45560 53193 45569 53227
rect 45569 53193 45603 53227
rect 45603 53193 45612 53227
rect 45560 53184 45612 53193
rect 47952 53184 48004 53236
rect 39488 53091 39540 53100
rect 39488 53057 39497 53091
rect 39497 53057 39531 53091
rect 39531 53057 39540 53091
rect 39488 53048 39540 53057
rect 42892 53116 42944 53168
rect 43352 53159 43404 53168
rect 43352 53125 43361 53159
rect 43361 53125 43395 53159
rect 43395 53125 43404 53159
rect 43352 53116 43404 53125
rect 37832 52980 37884 53032
rect 41420 52980 41472 53032
rect 41604 53048 41656 53100
rect 42616 53091 42668 53100
rect 42616 53057 42625 53091
rect 42625 53057 42659 53091
rect 42659 53057 42668 53091
rect 42616 53048 42668 53057
rect 42708 53091 42760 53100
rect 42708 53057 42717 53091
rect 42717 53057 42751 53091
rect 42751 53057 42760 53091
rect 42708 53048 42760 53057
rect 44180 53048 44232 53100
rect 46388 53116 46440 53168
rect 46940 53116 46992 53168
rect 50160 53184 50212 53236
rect 50620 53184 50672 53236
rect 45652 53091 45704 53100
rect 45652 53057 45661 53091
rect 45661 53057 45695 53091
rect 45695 53057 45704 53091
rect 45652 53048 45704 53057
rect 46204 53048 46256 53100
rect 47860 53091 47912 53100
rect 46112 52980 46164 53032
rect 47860 53057 47869 53091
rect 47869 53057 47903 53091
rect 47903 53057 47912 53091
rect 47860 53048 47912 53057
rect 48228 53091 48280 53100
rect 35532 52912 35584 52964
rect 41604 52912 41656 52964
rect 35716 52844 35768 52896
rect 48228 53057 48237 53091
rect 48237 53057 48271 53091
rect 48271 53057 48280 53091
rect 48228 53048 48280 53057
rect 48504 53048 48556 53100
rect 49884 53091 49936 53100
rect 49884 53057 49893 53091
rect 49893 53057 49927 53091
rect 49927 53057 49936 53091
rect 49884 53048 49936 53057
rect 50068 53091 50120 53100
rect 50068 53057 50077 53091
rect 50077 53057 50111 53091
rect 50111 53057 50120 53091
rect 50068 53048 50120 53057
rect 50712 53091 50764 53100
rect 50712 53057 50721 53091
rect 50721 53057 50755 53091
rect 50755 53057 50764 53091
rect 50712 53048 50764 53057
rect 48228 52912 48280 52964
rect 46296 52844 46348 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 65654 52742 65706 52794
rect 65718 52742 65770 52794
rect 65782 52742 65834 52794
rect 65846 52742 65898 52794
rect 65910 52742 65962 52794
rect 14096 52683 14148 52692
rect 14096 52649 14105 52683
rect 14105 52649 14139 52683
rect 14139 52649 14148 52683
rect 14096 52640 14148 52649
rect 15292 52640 15344 52692
rect 1400 52547 1452 52556
rect 1400 52513 1409 52547
rect 1409 52513 1443 52547
rect 1443 52513 1452 52547
rect 1400 52504 1452 52513
rect 1860 52547 1912 52556
rect 1860 52513 1869 52547
rect 1869 52513 1903 52547
rect 1903 52513 1912 52547
rect 1860 52504 1912 52513
rect 16580 52504 16632 52556
rect 17592 52504 17644 52556
rect 19340 52547 19392 52556
rect 19340 52513 19349 52547
rect 19349 52513 19383 52547
rect 19383 52513 19392 52547
rect 19340 52504 19392 52513
rect 21732 52572 21784 52624
rect 14280 52479 14332 52488
rect 14280 52445 14289 52479
rect 14289 52445 14323 52479
rect 14323 52445 14332 52479
rect 14280 52436 14332 52445
rect 16764 52436 16816 52488
rect 17132 52436 17184 52488
rect 18052 52479 18104 52488
rect 18052 52445 18061 52479
rect 18061 52445 18095 52479
rect 18095 52445 18104 52479
rect 18052 52436 18104 52445
rect 18144 52479 18196 52488
rect 18144 52445 18153 52479
rect 18153 52445 18187 52479
rect 18187 52445 18196 52479
rect 18144 52436 18196 52445
rect 1584 52411 1636 52420
rect 1584 52377 1593 52411
rect 1593 52377 1627 52411
rect 1627 52377 1636 52411
rect 1584 52368 1636 52377
rect 3516 52368 3568 52420
rect 16028 52411 16080 52420
rect 16028 52377 16037 52411
rect 16037 52377 16071 52411
rect 16071 52377 16080 52411
rect 16028 52368 16080 52377
rect 16304 52368 16356 52420
rect 18328 52368 18380 52420
rect 19432 52368 19484 52420
rect 21364 52411 21416 52420
rect 20720 52343 20772 52352
rect 20720 52309 20729 52343
rect 20729 52309 20763 52343
rect 20763 52309 20772 52343
rect 20720 52300 20772 52309
rect 21364 52377 21373 52411
rect 21373 52377 21407 52411
rect 21407 52377 21416 52411
rect 21364 52368 21416 52377
rect 21824 52479 21876 52488
rect 21824 52445 21838 52479
rect 21838 52445 21872 52479
rect 21872 52445 21876 52479
rect 21824 52436 21876 52445
rect 24400 52640 24452 52692
rect 28172 52683 28224 52692
rect 23664 52572 23716 52624
rect 24308 52572 24360 52624
rect 22468 52479 22520 52488
rect 22468 52445 22477 52479
rect 22477 52445 22511 52479
rect 22511 52445 22520 52479
rect 22468 52436 22520 52445
rect 23204 52436 23256 52488
rect 24216 52436 24268 52488
rect 24492 52479 24544 52488
rect 24492 52445 24501 52479
rect 24501 52445 24535 52479
rect 24535 52445 24544 52479
rect 24492 52436 24544 52445
rect 25412 52479 25464 52488
rect 25412 52445 25421 52479
rect 25421 52445 25455 52479
rect 25455 52445 25464 52479
rect 25412 52436 25464 52445
rect 26792 52479 26844 52488
rect 26792 52445 26801 52479
rect 26801 52445 26835 52479
rect 26835 52445 26844 52479
rect 26792 52436 26844 52445
rect 27436 52436 27488 52488
rect 28172 52649 28181 52683
rect 28181 52649 28215 52683
rect 28215 52649 28224 52683
rect 28172 52640 28224 52649
rect 28448 52640 28500 52692
rect 29092 52640 29144 52692
rect 29644 52640 29696 52692
rect 31392 52640 31444 52692
rect 33416 52640 33468 52692
rect 36636 52640 36688 52692
rect 43720 52683 43772 52692
rect 43720 52649 43729 52683
rect 43729 52649 43763 52683
rect 43763 52649 43772 52683
rect 43720 52640 43772 52649
rect 46204 52640 46256 52692
rect 48964 52640 49016 52692
rect 30564 52615 30616 52624
rect 30564 52581 30573 52615
rect 30573 52581 30607 52615
rect 30607 52581 30616 52615
rect 30564 52572 30616 52581
rect 35532 52572 35584 52624
rect 37280 52572 37332 52624
rect 37464 52572 37516 52624
rect 45744 52572 45796 52624
rect 28908 52436 28960 52488
rect 29552 52479 29604 52488
rect 29552 52445 29561 52479
rect 29561 52445 29595 52479
rect 29595 52445 29604 52479
rect 29552 52436 29604 52445
rect 30380 52479 30432 52488
rect 30380 52445 30389 52479
rect 30389 52445 30423 52479
rect 30423 52445 30432 52479
rect 30380 52436 30432 52445
rect 31116 52479 31168 52488
rect 31116 52445 31125 52479
rect 31125 52445 31159 52479
rect 31159 52445 31168 52479
rect 31116 52436 31168 52445
rect 31208 52436 31260 52488
rect 42616 52504 42668 52556
rect 45560 52504 45612 52556
rect 46112 52479 46164 52488
rect 46112 52445 46121 52479
rect 46121 52445 46155 52479
rect 46155 52445 46164 52479
rect 46112 52436 46164 52445
rect 46572 52436 46624 52488
rect 47584 52479 47636 52488
rect 47584 52445 47593 52479
rect 47593 52445 47627 52479
rect 47627 52445 47636 52479
rect 47584 52436 47636 52445
rect 50712 52436 50764 52488
rect 22560 52368 22612 52420
rect 23664 52368 23716 52420
rect 34152 52368 34204 52420
rect 35440 52411 35492 52420
rect 35440 52377 35449 52411
rect 35449 52377 35483 52411
rect 35483 52377 35492 52411
rect 35440 52368 35492 52377
rect 42340 52368 42392 52420
rect 43628 52368 43680 52420
rect 45468 52411 45520 52420
rect 45468 52377 45477 52411
rect 45477 52377 45511 52411
rect 45511 52377 45520 52411
rect 45468 52368 45520 52377
rect 45560 52368 45612 52420
rect 47860 52368 47912 52420
rect 24124 52300 24176 52352
rect 25136 52300 25188 52352
rect 28264 52300 28316 52352
rect 28908 52300 28960 52352
rect 32128 52300 32180 52352
rect 42892 52300 42944 52352
rect 44180 52343 44232 52352
rect 44180 52309 44189 52343
rect 44189 52309 44223 52343
rect 44223 52309 44232 52343
rect 44180 52300 44232 52309
rect 46940 52300 46992 52352
rect 47584 52300 47636 52352
rect 49792 52300 49844 52352
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 1584 52096 1636 52148
rect 2044 51960 2096 52012
rect 15016 51960 15068 52012
rect 18328 52003 18380 52012
rect 18328 51969 18337 52003
rect 18337 51969 18371 52003
rect 18371 51969 18380 52003
rect 18328 51960 18380 51969
rect 14372 51935 14424 51944
rect 14372 51901 14381 51935
rect 14381 51901 14415 51935
rect 14415 51901 14424 51935
rect 14372 51892 14424 51901
rect 17960 51824 18012 51876
rect 15752 51799 15804 51808
rect 15752 51765 15761 51799
rect 15761 51765 15795 51799
rect 15795 51765 15804 51799
rect 15752 51756 15804 51765
rect 17868 51756 17920 51808
rect 18420 51935 18472 51944
rect 18420 51901 18454 51935
rect 18454 51901 18472 51935
rect 18420 51892 18472 51901
rect 18604 51935 18656 51944
rect 18604 51901 18613 51935
rect 18613 51901 18647 51935
rect 18647 51901 18656 51935
rect 18604 51892 18656 51901
rect 18972 51892 19024 51944
rect 20076 52028 20128 52080
rect 20352 52028 20404 52080
rect 21364 52028 21416 52080
rect 23664 52071 23716 52080
rect 20720 51960 20772 52012
rect 23664 52037 23673 52071
rect 23673 52037 23707 52071
rect 23707 52037 23716 52071
rect 23664 52028 23716 52037
rect 29276 52028 29328 52080
rect 29552 52028 29604 52080
rect 32128 52071 32180 52080
rect 32128 52037 32137 52071
rect 32137 52037 32171 52071
rect 32171 52037 32180 52071
rect 32128 52028 32180 52037
rect 24308 52003 24360 52012
rect 20168 51892 20220 51944
rect 19248 51756 19300 51808
rect 19892 51799 19944 51808
rect 19892 51765 19901 51799
rect 19901 51765 19935 51799
rect 19935 51765 19944 51799
rect 19892 51756 19944 51765
rect 20076 51799 20128 51808
rect 20076 51765 20085 51799
rect 20085 51765 20119 51799
rect 20119 51765 20128 51799
rect 20076 51756 20128 51765
rect 22192 51756 22244 51808
rect 22468 51756 22520 51808
rect 22560 51756 22612 51808
rect 22928 51756 22980 51808
rect 24308 51969 24317 52003
rect 24317 51969 24351 52003
rect 24351 51969 24360 52003
rect 24308 51960 24360 51969
rect 24860 51960 24912 52012
rect 24584 51892 24636 51944
rect 24032 51824 24084 51876
rect 25320 51960 25372 52012
rect 25504 51960 25556 52012
rect 28080 52003 28132 52012
rect 28080 51969 28089 52003
rect 28089 51969 28123 52003
rect 28123 51969 28132 52003
rect 28080 51960 28132 51969
rect 28264 51960 28316 52012
rect 29736 51960 29788 52012
rect 34796 52028 34848 52080
rect 35992 52028 36044 52080
rect 42800 52028 42852 52080
rect 37556 51960 37608 52012
rect 37924 51960 37976 52012
rect 41236 52003 41288 52012
rect 41236 51969 41245 52003
rect 41245 51969 41279 52003
rect 41279 51969 41288 52003
rect 41236 51960 41288 51969
rect 41604 52003 41656 52012
rect 41604 51969 41613 52003
rect 41613 51969 41647 52003
rect 41647 51969 41656 52003
rect 41604 51960 41656 51969
rect 27804 51892 27856 51944
rect 28908 51892 28960 51944
rect 29368 51935 29420 51944
rect 29368 51901 29377 51935
rect 29377 51901 29411 51935
rect 29411 51901 29420 51935
rect 29368 51892 29420 51901
rect 25504 51824 25556 51876
rect 41696 51935 41748 51944
rect 41696 51901 41730 51935
rect 41730 51901 41748 51935
rect 43352 51960 43404 52012
rect 43720 52003 43772 52012
rect 43720 51969 43729 52003
rect 43729 51969 43763 52003
rect 43763 51969 43772 52003
rect 43720 51960 43772 51969
rect 45652 51960 45704 52012
rect 41696 51892 41748 51901
rect 24124 51756 24176 51808
rect 24768 51756 24820 51808
rect 31208 51824 31260 51876
rect 32496 51867 32548 51876
rect 32496 51833 32505 51867
rect 32505 51833 32539 51867
rect 32539 51833 32548 51867
rect 32496 51824 32548 51833
rect 35532 51867 35584 51876
rect 35532 51833 35541 51867
rect 35541 51833 35575 51867
rect 35575 51833 35584 51867
rect 35532 51824 35584 51833
rect 27804 51756 27856 51808
rect 30012 51756 30064 51808
rect 35624 51756 35676 51808
rect 37648 51756 37700 51808
rect 41604 51824 41656 51876
rect 41880 51867 41932 51876
rect 41880 51833 41889 51867
rect 41889 51833 41923 51867
rect 41923 51833 41932 51867
rect 41880 51824 41932 51833
rect 41236 51756 41288 51808
rect 43996 51892 44048 51944
rect 44088 51892 44140 51944
rect 46296 52003 46348 52012
rect 46296 51969 46305 52003
rect 46305 51969 46339 52003
rect 46339 51969 46348 52003
rect 46480 52003 46532 52012
rect 46296 51960 46348 51969
rect 46480 51969 46489 52003
rect 46489 51969 46523 52003
rect 46523 51969 46532 52003
rect 46480 51960 46532 51969
rect 47584 52003 47636 52012
rect 47584 51969 47593 52003
rect 47593 51969 47627 52003
rect 47627 51969 47636 52003
rect 47584 51960 47636 51969
rect 49792 52003 49844 52012
rect 49792 51969 49801 52003
rect 49801 51969 49835 52003
rect 49835 51969 49844 52003
rect 49792 51960 49844 51969
rect 51080 51960 51132 52012
rect 42892 51799 42944 51808
rect 42892 51765 42901 51799
rect 42901 51765 42935 51799
rect 42935 51765 42944 51799
rect 42892 51756 42944 51765
rect 46296 51824 46348 51876
rect 48964 51867 49016 51876
rect 48964 51833 48973 51867
rect 48973 51833 49007 51867
rect 49007 51833 49016 51867
rect 48964 51824 49016 51833
rect 48228 51756 48280 51808
rect 50528 51756 50580 51808
rect 66076 51756 66128 51808
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 65654 51654 65706 51706
rect 65718 51654 65770 51706
rect 65782 51654 65834 51706
rect 65846 51654 65898 51706
rect 65910 51654 65962 51706
rect 15016 51595 15068 51604
rect 15016 51561 15025 51595
rect 15025 51561 15059 51595
rect 15059 51561 15068 51595
rect 15016 51552 15068 51561
rect 18052 51552 18104 51604
rect 19432 51552 19484 51604
rect 26792 51595 26844 51604
rect 26792 51561 26801 51595
rect 26801 51561 26835 51595
rect 26835 51561 26844 51595
rect 26792 51552 26844 51561
rect 17960 51484 18012 51536
rect 19248 51484 19300 51536
rect 21824 51484 21876 51536
rect 26332 51484 26384 51536
rect 18144 51416 18196 51468
rect 24768 51416 24820 51468
rect 28080 51416 28132 51468
rect 29644 51416 29696 51468
rect 34888 51484 34940 51536
rect 35992 51527 36044 51536
rect 35992 51493 36001 51527
rect 36001 51493 36035 51527
rect 36035 51493 36044 51527
rect 35992 51484 36044 51493
rect 36452 51527 36504 51536
rect 36452 51493 36461 51527
rect 36461 51493 36495 51527
rect 36495 51493 36504 51527
rect 36452 51484 36504 51493
rect 37924 51552 37976 51604
rect 41696 51552 41748 51604
rect 30748 51459 30800 51468
rect 30748 51425 30757 51459
rect 30757 51425 30791 51459
rect 30791 51425 30800 51459
rect 30748 51416 30800 51425
rect 34428 51416 34480 51468
rect 15752 51391 15804 51400
rect 15752 51357 15761 51391
rect 15761 51357 15795 51391
rect 15795 51357 15804 51391
rect 15752 51348 15804 51357
rect 16580 51348 16632 51400
rect 16764 51391 16816 51400
rect 16764 51357 16773 51391
rect 16773 51357 16807 51391
rect 16807 51357 16816 51391
rect 16764 51348 16816 51357
rect 18420 51348 18472 51400
rect 20076 51348 20128 51400
rect 20352 51348 20404 51400
rect 25136 51391 25188 51400
rect 25136 51357 25170 51391
rect 25170 51357 25188 51391
rect 17408 51280 17460 51332
rect 20536 51323 20588 51332
rect 20536 51289 20545 51323
rect 20545 51289 20579 51323
rect 20579 51289 20588 51323
rect 20536 51280 20588 51289
rect 25136 51348 25188 51357
rect 26240 51348 26292 51400
rect 27988 51391 28040 51400
rect 27988 51357 27997 51391
rect 27997 51357 28031 51391
rect 28031 51357 28040 51391
rect 27988 51348 28040 51357
rect 28264 51391 28316 51400
rect 28264 51357 28273 51391
rect 28273 51357 28307 51391
rect 28307 51357 28316 51391
rect 28264 51348 28316 51357
rect 24952 51280 25004 51332
rect 13820 51212 13872 51264
rect 14648 51212 14700 51264
rect 14740 51212 14792 51264
rect 24400 51212 24452 51264
rect 30472 51391 30524 51400
rect 30472 51357 30481 51391
rect 30481 51357 30515 51391
rect 30515 51357 30524 51391
rect 30472 51348 30524 51357
rect 32036 51348 32088 51400
rect 32772 51391 32824 51400
rect 32772 51357 32781 51391
rect 32781 51357 32815 51391
rect 32815 51357 32824 51391
rect 32772 51348 32824 51357
rect 34704 51391 34756 51400
rect 34704 51357 34713 51391
rect 34713 51357 34747 51391
rect 34747 51357 34756 51391
rect 34704 51348 34756 51357
rect 34888 51391 34940 51400
rect 34888 51357 34897 51391
rect 34897 51357 34931 51391
rect 34931 51357 34940 51391
rect 34888 51348 34940 51357
rect 35624 51348 35676 51400
rect 35808 51391 35860 51400
rect 35808 51357 35817 51391
rect 35817 51357 35851 51391
rect 35851 51357 35860 51391
rect 35808 51348 35860 51357
rect 36360 51348 36412 51400
rect 36728 51391 36780 51400
rect 36728 51357 36737 51391
rect 36737 51357 36771 51391
rect 36771 51357 36780 51391
rect 36728 51348 36780 51357
rect 37648 51391 37700 51400
rect 37648 51357 37657 51391
rect 37657 51357 37691 51391
rect 37691 51357 37700 51391
rect 37648 51348 37700 51357
rect 38660 51391 38712 51400
rect 32128 51280 32180 51332
rect 34152 51255 34204 51264
rect 34152 51221 34161 51255
rect 34161 51221 34195 51255
rect 34195 51221 34204 51255
rect 36084 51280 36136 51332
rect 37096 51280 37148 51332
rect 38660 51357 38669 51391
rect 38669 51357 38703 51391
rect 38703 51357 38712 51391
rect 38660 51348 38712 51357
rect 38844 51391 38896 51400
rect 38844 51357 38853 51391
rect 38853 51357 38887 51391
rect 38887 51357 38896 51391
rect 38844 51348 38896 51357
rect 41604 51484 41656 51536
rect 51080 51527 51132 51536
rect 42524 51459 42576 51468
rect 42524 51425 42533 51459
rect 42533 51425 42567 51459
rect 42567 51425 42576 51459
rect 42524 51416 42576 51425
rect 51080 51493 51089 51527
rect 51089 51493 51123 51527
rect 51123 51493 51132 51527
rect 51080 51484 51132 51493
rect 43904 51416 43956 51468
rect 50068 51416 50120 51468
rect 50528 51416 50580 51468
rect 42340 51391 42392 51400
rect 42340 51357 42349 51391
rect 42349 51357 42383 51391
rect 42383 51357 42392 51391
rect 42340 51348 42392 51357
rect 42616 51391 42668 51400
rect 42616 51357 42625 51391
rect 42625 51357 42659 51391
rect 42659 51357 42668 51391
rect 42616 51348 42668 51357
rect 42984 51391 43036 51400
rect 42984 51357 42993 51391
rect 42993 51357 43027 51391
rect 43027 51357 43036 51391
rect 42984 51348 43036 51357
rect 43628 51348 43680 51400
rect 43812 51391 43864 51400
rect 43812 51357 43821 51391
rect 43821 51357 43855 51391
rect 43855 51357 43864 51391
rect 43996 51391 44048 51400
rect 43812 51348 43864 51357
rect 43996 51357 44005 51391
rect 44005 51357 44039 51391
rect 44039 51357 44048 51391
rect 43996 51348 44048 51357
rect 44088 51391 44140 51400
rect 44088 51357 44097 51391
rect 44097 51357 44131 51391
rect 44131 51357 44140 51391
rect 44088 51348 44140 51357
rect 41880 51280 41932 51332
rect 45192 51391 45244 51400
rect 45192 51357 45201 51391
rect 45201 51357 45235 51391
rect 45235 51357 45244 51391
rect 45192 51348 45244 51357
rect 45468 51348 45520 51400
rect 46112 51348 46164 51400
rect 46572 51348 46624 51400
rect 48412 51348 48464 51400
rect 45652 51280 45704 51332
rect 50160 51280 50212 51332
rect 66444 51323 66496 51332
rect 66444 51289 66453 51323
rect 66453 51289 66487 51323
rect 66487 51289 66496 51323
rect 66444 51280 66496 51289
rect 68100 51323 68152 51332
rect 68100 51289 68109 51323
rect 68109 51289 68143 51323
rect 68143 51289 68152 51323
rect 68100 51280 68152 51289
rect 34152 51212 34204 51221
rect 35532 51212 35584 51264
rect 35716 51212 35768 51264
rect 38752 51212 38804 51264
rect 43168 51212 43220 51264
rect 43812 51212 43864 51264
rect 43904 51212 43956 51264
rect 45836 51212 45888 51264
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 14372 51008 14424 51060
rect 16764 51008 16816 51060
rect 17408 51051 17460 51060
rect 17408 51017 17417 51051
rect 17417 51017 17451 51051
rect 17451 51017 17460 51051
rect 17408 51008 17460 51017
rect 20444 51008 20496 51060
rect 23756 51008 23808 51060
rect 24032 51008 24084 51060
rect 25412 51008 25464 51060
rect 28080 51008 28132 51060
rect 30472 51008 30524 51060
rect 31392 51008 31444 51060
rect 14096 50872 14148 50924
rect 14648 50915 14700 50924
rect 14648 50881 14657 50915
rect 14657 50881 14691 50915
rect 14691 50881 14700 50915
rect 14648 50872 14700 50881
rect 16856 50915 16908 50924
rect 16856 50881 16865 50915
rect 16865 50881 16899 50915
rect 16899 50881 16908 50915
rect 16856 50872 16908 50881
rect 17316 50872 17368 50924
rect 17592 50915 17644 50924
rect 17592 50881 17601 50915
rect 17601 50881 17635 50915
rect 17635 50881 17644 50915
rect 17592 50872 17644 50881
rect 20260 50872 20312 50924
rect 20996 50915 21048 50924
rect 20996 50881 21005 50915
rect 21005 50881 21039 50915
rect 21039 50881 21048 50915
rect 20996 50872 21048 50881
rect 24400 50872 24452 50924
rect 24676 50872 24728 50924
rect 25044 50872 25096 50924
rect 26332 50940 26384 50992
rect 31116 50983 31168 50992
rect 25320 50804 25372 50856
rect 26240 50915 26292 50924
rect 26240 50881 26249 50915
rect 26249 50881 26283 50915
rect 26283 50881 26292 50915
rect 26240 50872 26292 50881
rect 27620 50872 27672 50924
rect 31116 50949 31125 50983
rect 31125 50949 31159 50983
rect 31159 50949 31168 50983
rect 31116 50940 31168 50949
rect 31208 50940 31260 50992
rect 34704 50940 34756 50992
rect 35440 50940 35492 50992
rect 35808 50940 35860 50992
rect 36820 51008 36872 51060
rect 46388 51051 46440 51060
rect 28908 50804 28960 50856
rect 30564 50872 30616 50924
rect 34152 50915 34204 50924
rect 34152 50881 34161 50915
rect 34161 50881 34195 50915
rect 34195 50881 34204 50915
rect 34152 50872 34204 50881
rect 34428 50847 34480 50856
rect 29552 50736 29604 50788
rect 14280 50668 14332 50720
rect 19524 50711 19576 50720
rect 19524 50677 19533 50711
rect 19533 50677 19567 50711
rect 19567 50677 19576 50711
rect 19524 50668 19576 50677
rect 31300 50668 31352 50720
rect 34428 50813 34437 50847
rect 34437 50813 34471 50847
rect 34471 50813 34480 50847
rect 34428 50804 34480 50813
rect 36544 50872 36596 50924
rect 46388 51017 46397 51051
rect 46397 51017 46431 51051
rect 46431 51017 46440 51051
rect 46388 51008 46440 51017
rect 46664 51008 46716 51060
rect 66444 51051 66496 51060
rect 66444 51017 66453 51051
rect 66453 51017 66487 51051
rect 66487 51017 66496 51051
rect 66444 51008 66496 51017
rect 38476 50872 38528 50924
rect 46296 50983 46348 50992
rect 46296 50949 46305 50983
rect 46305 50949 46339 50983
rect 46339 50949 46348 50983
rect 46296 50940 46348 50949
rect 39488 50915 39540 50924
rect 39488 50881 39497 50915
rect 39497 50881 39531 50915
rect 39531 50881 39540 50915
rect 39488 50872 39540 50881
rect 41052 50872 41104 50924
rect 43628 50872 43680 50924
rect 43904 50915 43956 50924
rect 43904 50881 43913 50915
rect 43913 50881 43947 50915
rect 43947 50881 43956 50915
rect 43904 50872 43956 50881
rect 44088 50872 44140 50924
rect 45652 50872 45704 50924
rect 47676 50915 47728 50924
rect 47676 50881 47685 50915
rect 47685 50881 47719 50915
rect 47719 50881 47728 50915
rect 47676 50872 47728 50881
rect 48228 50872 48280 50924
rect 34244 50779 34296 50788
rect 34244 50745 34253 50779
rect 34253 50745 34287 50779
rect 34287 50745 34296 50779
rect 34244 50736 34296 50745
rect 36636 50779 36688 50788
rect 36636 50745 36645 50779
rect 36645 50745 36679 50779
rect 36679 50745 36688 50779
rect 36636 50736 36688 50745
rect 35716 50711 35768 50720
rect 35716 50677 35725 50711
rect 35725 50677 35759 50711
rect 35759 50677 35768 50711
rect 42800 50804 42852 50856
rect 43996 50847 44048 50856
rect 43996 50813 44005 50847
rect 44005 50813 44039 50847
rect 44039 50813 44048 50847
rect 43996 50804 44048 50813
rect 38016 50779 38068 50788
rect 38016 50745 38025 50779
rect 38025 50745 38059 50779
rect 38059 50745 38068 50779
rect 38016 50736 38068 50745
rect 38752 50736 38804 50788
rect 41604 50779 41656 50788
rect 41604 50745 41613 50779
rect 41613 50745 41647 50779
rect 41647 50745 41656 50779
rect 41604 50736 41656 50745
rect 42616 50736 42668 50788
rect 47032 50804 47084 50856
rect 48412 50804 48464 50856
rect 50160 50915 50212 50924
rect 50160 50881 50169 50915
rect 50169 50881 50203 50915
rect 50203 50881 50212 50915
rect 50160 50872 50212 50881
rect 51540 50872 51592 50924
rect 66812 50872 66864 50924
rect 48780 50847 48832 50856
rect 48780 50813 48789 50847
rect 48789 50813 48823 50847
rect 48823 50813 48832 50847
rect 48780 50804 48832 50813
rect 50988 50804 51040 50856
rect 46204 50736 46256 50788
rect 47124 50736 47176 50788
rect 35716 50668 35768 50677
rect 43444 50668 43496 50720
rect 47308 50668 47360 50720
rect 48596 50711 48648 50720
rect 48596 50677 48605 50711
rect 48605 50677 48639 50711
rect 48639 50677 48648 50711
rect 48596 50668 48648 50677
rect 49056 50711 49108 50720
rect 49056 50677 49065 50711
rect 49065 50677 49099 50711
rect 49099 50677 49108 50711
rect 49056 50668 49108 50677
rect 52736 50711 52788 50720
rect 52736 50677 52745 50711
rect 52745 50677 52779 50711
rect 52779 50677 52788 50711
rect 52736 50668 52788 50677
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 65654 50566 65706 50618
rect 65718 50566 65770 50618
rect 65782 50566 65834 50618
rect 65846 50566 65898 50618
rect 65910 50566 65962 50618
rect 24400 50464 24452 50516
rect 27620 50507 27672 50516
rect 20996 50396 21048 50448
rect 27620 50473 27629 50507
rect 27629 50473 27663 50507
rect 27663 50473 27672 50507
rect 27620 50464 27672 50473
rect 32496 50507 32548 50516
rect 32496 50473 32505 50507
rect 32505 50473 32539 50507
rect 32539 50473 32548 50507
rect 32496 50464 32548 50473
rect 36820 50464 36872 50516
rect 37096 50464 37148 50516
rect 21456 50328 21508 50380
rect 14096 50260 14148 50312
rect 15108 50303 15160 50312
rect 15108 50269 15117 50303
rect 15117 50269 15151 50303
rect 15151 50269 15160 50303
rect 15108 50260 15160 50269
rect 15200 50303 15252 50312
rect 15200 50269 15209 50303
rect 15209 50269 15243 50303
rect 15243 50269 15252 50303
rect 15200 50260 15252 50269
rect 18512 50260 18564 50312
rect 19340 50260 19392 50312
rect 19524 50303 19576 50312
rect 19524 50269 19558 50303
rect 19558 50269 19576 50303
rect 19524 50260 19576 50269
rect 20076 50260 20128 50312
rect 22560 50260 22612 50312
rect 24124 50328 24176 50380
rect 29736 50396 29788 50448
rect 13820 50192 13872 50244
rect 18604 50192 18656 50244
rect 12440 50124 12492 50176
rect 15384 50167 15436 50176
rect 15384 50133 15393 50167
rect 15393 50133 15427 50167
rect 15427 50133 15436 50167
rect 15384 50124 15436 50133
rect 16580 50124 16632 50176
rect 17684 50124 17736 50176
rect 22284 50192 22336 50244
rect 23020 50303 23072 50312
rect 23020 50269 23029 50303
rect 23029 50269 23063 50303
rect 23063 50269 23072 50303
rect 23020 50260 23072 50269
rect 23388 50260 23440 50312
rect 23480 50260 23532 50312
rect 24032 50260 24084 50312
rect 27804 50303 27856 50312
rect 27804 50269 27813 50303
rect 27813 50269 27847 50303
rect 27847 50269 27856 50303
rect 27804 50260 27856 50269
rect 27988 50328 28040 50380
rect 37648 50396 37700 50448
rect 38476 50464 38528 50516
rect 40500 50464 40552 50516
rect 41052 50507 41104 50516
rect 41052 50473 41061 50507
rect 41061 50473 41095 50507
rect 41095 50473 41104 50507
rect 41052 50464 41104 50473
rect 41788 50464 41840 50516
rect 47032 50464 47084 50516
rect 47308 50507 47360 50516
rect 47308 50473 47317 50507
rect 47317 50473 47351 50507
rect 47351 50473 47360 50507
rect 47308 50464 47360 50473
rect 43444 50396 43496 50448
rect 49056 50464 49108 50516
rect 50068 50464 50120 50516
rect 50988 50464 51040 50516
rect 29920 50303 29972 50312
rect 29920 50269 29929 50303
rect 29929 50269 29963 50303
rect 29963 50269 29972 50303
rect 29920 50260 29972 50269
rect 30012 50260 30064 50312
rect 30288 50260 30340 50312
rect 32588 50260 32640 50312
rect 19984 50124 20036 50176
rect 22376 50167 22428 50176
rect 22376 50133 22385 50167
rect 22385 50133 22419 50167
rect 22419 50133 22428 50167
rect 22376 50124 22428 50133
rect 25872 50192 25924 50244
rect 36084 50303 36136 50312
rect 36084 50269 36093 50303
rect 36093 50269 36127 50303
rect 36127 50269 36136 50303
rect 36084 50260 36136 50269
rect 36544 50260 36596 50312
rect 38568 50303 38620 50312
rect 38568 50269 38577 50303
rect 38577 50269 38611 50303
rect 38611 50269 38620 50303
rect 38568 50260 38620 50269
rect 41604 50328 41656 50380
rect 39672 50260 39724 50312
rect 41328 50260 41380 50312
rect 41880 50260 41932 50312
rect 42432 50260 42484 50312
rect 45836 50303 45888 50312
rect 45836 50269 45845 50303
rect 45845 50269 45879 50303
rect 45879 50269 45888 50303
rect 45836 50260 45888 50269
rect 46296 50260 46348 50312
rect 47124 50371 47176 50380
rect 47124 50337 47133 50371
rect 47133 50337 47167 50371
rect 47167 50337 47176 50371
rect 47124 50328 47176 50337
rect 34428 50192 34480 50244
rect 36636 50192 36688 50244
rect 37556 50235 37608 50244
rect 37556 50201 37565 50235
rect 37565 50201 37599 50235
rect 37599 50201 37608 50235
rect 37556 50192 37608 50201
rect 29920 50124 29972 50176
rect 33324 50124 33376 50176
rect 35716 50124 35768 50176
rect 37096 50124 37148 50176
rect 37464 50124 37516 50176
rect 37740 50124 37792 50176
rect 38016 50124 38068 50176
rect 44088 50192 44140 50244
rect 45652 50192 45704 50244
rect 47768 50260 47820 50312
rect 48780 50396 48832 50448
rect 48228 50328 48280 50380
rect 48320 50192 48372 50244
rect 48596 50260 48648 50312
rect 50160 50260 50212 50312
rect 50620 50260 50672 50312
rect 51356 50260 51408 50312
rect 52736 50260 52788 50312
rect 49792 50192 49844 50244
rect 41972 50124 42024 50176
rect 43076 50124 43128 50176
rect 45928 50167 45980 50176
rect 45928 50133 45937 50167
rect 45937 50133 45971 50167
rect 45971 50133 45980 50167
rect 45928 50124 45980 50133
rect 46112 50124 46164 50176
rect 47492 50167 47544 50176
rect 47492 50133 47501 50167
rect 47501 50133 47535 50167
rect 47535 50133 47544 50167
rect 47492 50124 47544 50133
rect 48136 50167 48188 50176
rect 48136 50133 48145 50167
rect 48145 50133 48179 50167
rect 48179 50133 48188 50167
rect 48136 50124 48188 50133
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 3516 49920 3568 49972
rect 17684 49920 17736 49972
rect 12440 49827 12492 49836
rect 12440 49793 12449 49827
rect 12449 49793 12483 49827
rect 12483 49793 12492 49827
rect 12440 49784 12492 49793
rect 12992 49784 13044 49836
rect 14280 49827 14332 49836
rect 14280 49793 14289 49827
rect 14289 49793 14323 49827
rect 14323 49793 14332 49827
rect 14280 49784 14332 49793
rect 14372 49784 14424 49836
rect 15108 49784 15160 49836
rect 16856 49827 16908 49836
rect 16856 49793 16865 49827
rect 16865 49793 16899 49827
rect 16899 49793 16908 49827
rect 16856 49784 16908 49793
rect 13820 49691 13872 49700
rect 13820 49657 13829 49691
rect 13829 49657 13863 49691
rect 13863 49657 13872 49691
rect 13820 49648 13872 49657
rect 17592 49759 17644 49768
rect 17592 49725 17601 49759
rect 17601 49725 17635 49759
rect 17635 49725 17644 49759
rect 19984 49920 20036 49972
rect 20260 49963 20312 49972
rect 20260 49929 20269 49963
rect 20269 49929 20303 49963
rect 20303 49929 20312 49963
rect 20260 49920 20312 49929
rect 24952 49963 25004 49972
rect 24952 49929 24961 49963
rect 24961 49929 24995 49963
rect 24995 49929 25004 49963
rect 24952 49920 25004 49929
rect 25136 49920 25188 49972
rect 25504 49920 25556 49972
rect 18604 49827 18656 49836
rect 18604 49793 18638 49827
rect 18638 49793 18656 49827
rect 22284 49852 22336 49904
rect 18604 49784 18656 49793
rect 20260 49784 20312 49836
rect 17592 49716 17644 49725
rect 18972 49716 19024 49768
rect 20628 49716 20680 49768
rect 18236 49691 18288 49700
rect 18236 49657 18245 49691
rect 18245 49657 18279 49691
rect 18279 49657 18288 49691
rect 18236 49648 18288 49657
rect 22836 49716 22888 49768
rect 24400 49784 24452 49836
rect 27344 49784 27396 49836
rect 29184 49784 29236 49836
rect 22560 49648 22612 49700
rect 23020 49648 23072 49700
rect 16856 49623 16908 49632
rect 16856 49589 16865 49623
rect 16865 49589 16899 49623
rect 16899 49589 16908 49623
rect 16856 49580 16908 49589
rect 20076 49623 20128 49632
rect 20076 49589 20085 49623
rect 20085 49589 20119 49623
rect 20119 49589 20128 49623
rect 20076 49580 20128 49589
rect 26056 49623 26108 49632
rect 26056 49589 26065 49623
rect 26065 49589 26099 49623
rect 26099 49589 26108 49623
rect 26056 49580 26108 49589
rect 28632 49623 28684 49632
rect 28632 49589 28641 49623
rect 28641 49589 28675 49623
rect 28675 49589 28684 49623
rect 28632 49580 28684 49589
rect 32588 49920 32640 49972
rect 37372 49920 37424 49972
rect 37648 49920 37700 49972
rect 30104 49784 30156 49836
rect 36084 49852 36136 49904
rect 30932 49784 30984 49836
rect 32036 49784 32088 49836
rect 34244 49827 34296 49836
rect 29736 49716 29788 49768
rect 31392 49716 31444 49768
rect 34244 49793 34253 49827
rect 34253 49793 34287 49827
rect 34287 49793 34296 49827
rect 34244 49784 34296 49793
rect 35440 49827 35492 49836
rect 35440 49793 35449 49827
rect 35449 49793 35483 49827
rect 35483 49793 35492 49827
rect 35440 49784 35492 49793
rect 35532 49784 35584 49836
rect 35808 49784 35860 49836
rect 36544 49827 36596 49836
rect 36544 49793 36553 49827
rect 36553 49793 36587 49827
rect 36587 49793 36596 49827
rect 36544 49784 36596 49793
rect 37556 49852 37608 49904
rect 38292 49895 38344 49904
rect 38292 49861 38301 49895
rect 38301 49861 38335 49895
rect 38335 49861 38344 49895
rect 38292 49852 38344 49861
rect 41696 49895 41748 49904
rect 36452 49716 36504 49768
rect 37096 49716 37148 49768
rect 39672 49784 39724 49836
rect 41696 49861 41722 49895
rect 41722 49861 41748 49895
rect 41696 49852 41748 49861
rect 45928 49920 45980 49972
rect 43444 49852 43496 49904
rect 44640 49852 44692 49904
rect 46388 49920 46440 49972
rect 49332 49920 49384 49972
rect 51356 49963 51408 49972
rect 51356 49929 51365 49963
rect 51365 49929 51399 49963
rect 51399 49929 51408 49963
rect 51356 49920 51408 49929
rect 42432 49827 42484 49836
rect 42432 49793 42441 49827
rect 42441 49793 42475 49827
rect 42475 49793 42484 49827
rect 42432 49784 42484 49793
rect 44916 49827 44968 49836
rect 33508 49580 33560 49632
rect 34796 49623 34848 49632
rect 34796 49589 34805 49623
rect 34805 49589 34839 49623
rect 34839 49589 34848 49623
rect 34796 49580 34848 49589
rect 37280 49580 37332 49632
rect 44180 49648 44232 49700
rect 44916 49793 44925 49827
rect 44925 49793 44959 49827
rect 44959 49793 44968 49827
rect 44916 49784 44968 49793
rect 45008 49827 45060 49836
rect 47676 49852 47728 49904
rect 45008 49793 45043 49827
rect 45043 49793 45060 49827
rect 45008 49784 45060 49793
rect 45652 49716 45704 49768
rect 46296 49716 46348 49768
rect 47768 49759 47820 49768
rect 47768 49725 47777 49759
rect 47777 49725 47811 49759
rect 47811 49725 47820 49759
rect 47768 49716 47820 49725
rect 45100 49648 45152 49700
rect 49332 49784 49384 49836
rect 50620 49784 50672 49836
rect 51356 49784 51408 49836
rect 52092 49827 52144 49836
rect 52092 49793 52101 49827
rect 52101 49793 52135 49827
rect 52135 49793 52144 49827
rect 52092 49784 52144 49793
rect 42064 49580 42116 49632
rect 42616 49623 42668 49632
rect 42616 49589 42625 49623
rect 42625 49589 42659 49623
rect 42659 49589 42668 49623
rect 42616 49580 42668 49589
rect 43536 49623 43588 49632
rect 43536 49589 43545 49623
rect 43545 49589 43579 49623
rect 43579 49589 43588 49623
rect 43536 49580 43588 49589
rect 44916 49580 44968 49632
rect 45376 49580 45428 49632
rect 46480 49580 46532 49632
rect 48228 49580 48280 49632
rect 50252 49759 50304 49768
rect 50252 49725 50261 49759
rect 50261 49725 50295 49759
rect 50295 49725 50304 49759
rect 50252 49716 50304 49725
rect 49056 49580 49108 49632
rect 50068 49623 50120 49632
rect 50068 49589 50077 49623
rect 50077 49589 50111 49623
rect 50111 49589 50120 49623
rect 50068 49580 50120 49589
rect 52000 49580 52052 49632
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 65654 49478 65706 49530
rect 65718 49478 65770 49530
rect 65782 49478 65834 49530
rect 65846 49478 65898 49530
rect 65910 49478 65962 49530
rect 14372 49419 14424 49428
rect 14372 49385 14381 49419
rect 14381 49385 14415 49419
rect 14415 49385 14424 49419
rect 14372 49376 14424 49385
rect 17592 49376 17644 49428
rect 18512 49419 18564 49428
rect 13820 49240 13872 49292
rect 13268 49215 13320 49224
rect 13268 49181 13277 49215
rect 13277 49181 13311 49215
rect 13311 49181 13320 49215
rect 13268 49172 13320 49181
rect 15384 49240 15436 49292
rect 18512 49385 18521 49419
rect 18521 49385 18555 49419
rect 18555 49385 18564 49419
rect 18512 49376 18564 49385
rect 19340 49419 19392 49428
rect 19340 49385 19349 49419
rect 19349 49385 19383 49419
rect 19383 49385 19392 49419
rect 19340 49376 19392 49385
rect 23020 49419 23072 49428
rect 23020 49385 23029 49419
rect 23029 49385 23063 49419
rect 23063 49385 23072 49419
rect 23020 49376 23072 49385
rect 30932 49376 30984 49428
rect 28724 49308 28776 49360
rect 15200 49172 15252 49224
rect 16856 49172 16908 49224
rect 17316 49172 17368 49224
rect 35440 49376 35492 49428
rect 40040 49376 40092 49428
rect 41328 49376 41380 49428
rect 43536 49376 43588 49428
rect 46296 49419 46348 49428
rect 40132 49351 40184 49360
rect 16028 49104 16080 49156
rect 16580 49147 16632 49156
rect 16580 49113 16614 49147
rect 16614 49113 16632 49147
rect 20536 49172 20588 49224
rect 22192 49172 22244 49224
rect 23296 49172 23348 49224
rect 24860 49215 24912 49224
rect 24860 49181 24869 49215
rect 24869 49181 24903 49215
rect 24903 49181 24912 49215
rect 24860 49172 24912 49181
rect 26056 49172 26108 49224
rect 26332 49172 26384 49224
rect 28632 49172 28684 49224
rect 30288 49215 30340 49224
rect 30288 49181 30297 49215
rect 30297 49181 30331 49215
rect 30331 49181 30340 49215
rect 30288 49172 30340 49181
rect 31300 49215 31352 49224
rect 31300 49181 31309 49215
rect 31309 49181 31343 49215
rect 31343 49181 31352 49215
rect 31300 49172 31352 49181
rect 32588 49215 32640 49224
rect 32588 49181 32597 49215
rect 32597 49181 32631 49215
rect 32631 49181 32640 49215
rect 32588 49172 32640 49181
rect 34704 49215 34756 49224
rect 34704 49181 34713 49215
rect 34713 49181 34747 49215
rect 34747 49181 34756 49215
rect 34704 49172 34756 49181
rect 36636 49172 36688 49224
rect 16580 49104 16632 49113
rect 20260 49104 20312 49156
rect 22376 49104 22428 49156
rect 30840 49104 30892 49156
rect 32680 49104 32732 49156
rect 33048 49104 33100 49156
rect 33416 49104 33468 49156
rect 34612 49104 34664 49156
rect 36544 49104 36596 49156
rect 37648 49104 37700 49156
rect 13176 49036 13228 49088
rect 23296 49036 23348 49088
rect 27620 49036 27672 49088
rect 29092 49036 29144 49088
rect 33508 49036 33560 49088
rect 37280 49079 37332 49088
rect 37280 49045 37289 49079
rect 37289 49045 37323 49079
rect 37323 49045 37332 49079
rect 37280 49036 37332 49045
rect 37464 49036 37516 49088
rect 38292 49215 38344 49224
rect 38292 49181 38301 49215
rect 38301 49181 38335 49215
rect 38335 49181 38344 49215
rect 38292 49172 38344 49181
rect 39672 49172 39724 49224
rect 40132 49317 40141 49351
rect 40141 49317 40175 49351
rect 40175 49317 40184 49351
rect 40132 49308 40184 49317
rect 41696 49308 41748 49360
rect 42616 49308 42668 49360
rect 41420 49215 41472 49224
rect 41420 49181 41429 49215
rect 41429 49181 41463 49215
rect 41463 49181 41472 49215
rect 41420 49172 41472 49181
rect 41696 49172 41748 49224
rect 41972 49215 42024 49224
rect 41972 49181 41981 49215
rect 41981 49181 42015 49215
rect 42015 49181 42024 49215
rect 41972 49172 42024 49181
rect 43444 49215 43496 49224
rect 43444 49181 43453 49215
rect 43453 49181 43487 49215
rect 43487 49181 43496 49215
rect 43444 49172 43496 49181
rect 45560 49308 45612 49360
rect 46296 49385 46305 49419
rect 46305 49385 46339 49419
rect 46339 49385 46348 49419
rect 46296 49376 46348 49385
rect 48320 49376 48372 49428
rect 52092 49376 52144 49428
rect 47492 49308 47544 49360
rect 43904 49215 43956 49224
rect 43904 49181 43913 49215
rect 43913 49181 43947 49215
rect 43947 49181 43956 49215
rect 43904 49172 43956 49181
rect 45376 49215 45428 49224
rect 45376 49181 45385 49215
rect 45385 49181 45419 49215
rect 45419 49181 45428 49215
rect 45376 49172 45428 49181
rect 45652 49215 45704 49224
rect 45652 49181 45661 49215
rect 45661 49181 45695 49215
rect 45695 49181 45704 49215
rect 45652 49172 45704 49181
rect 46480 49215 46532 49224
rect 45100 49104 45152 49156
rect 46480 49181 46489 49215
rect 46489 49181 46523 49215
rect 46523 49181 46532 49215
rect 46480 49172 46532 49181
rect 47676 49172 47728 49224
rect 48596 49172 48648 49224
rect 49332 49215 49384 49224
rect 49332 49181 49341 49215
rect 49341 49181 49375 49215
rect 49375 49181 49384 49215
rect 49332 49172 49384 49181
rect 50252 49172 50304 49224
rect 40224 49036 40276 49088
rect 40316 49036 40368 49088
rect 45376 49036 45428 49088
rect 45928 49036 45980 49088
rect 51540 49172 51592 49224
rect 51632 49172 51684 49224
rect 52000 49215 52052 49224
rect 52000 49181 52034 49215
rect 52034 49181 52052 49215
rect 52000 49172 52052 49181
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 12992 48875 13044 48884
rect 12992 48841 13001 48875
rect 13001 48841 13035 48875
rect 13035 48841 13044 48875
rect 12992 48832 13044 48841
rect 20720 48832 20772 48884
rect 26332 48875 26384 48884
rect 13268 48764 13320 48816
rect 20812 48764 20864 48816
rect 26332 48841 26341 48875
rect 26341 48841 26375 48875
rect 26375 48841 26384 48875
rect 26332 48832 26384 48841
rect 27344 48875 27396 48884
rect 27344 48841 27353 48875
rect 27353 48841 27387 48875
rect 27387 48841 27396 48875
rect 27344 48832 27396 48841
rect 29184 48832 29236 48884
rect 34612 48875 34664 48884
rect 34612 48841 34621 48875
rect 34621 48841 34655 48875
rect 34655 48841 34664 48875
rect 34612 48832 34664 48841
rect 13176 48739 13228 48748
rect 13176 48705 13185 48739
rect 13185 48705 13219 48739
rect 13219 48705 13228 48739
rect 13176 48696 13228 48705
rect 17132 48739 17184 48748
rect 17132 48705 17141 48739
rect 17141 48705 17175 48739
rect 17175 48705 17184 48739
rect 17132 48696 17184 48705
rect 19984 48696 20036 48748
rect 20260 48739 20312 48748
rect 20260 48705 20269 48739
rect 20269 48705 20303 48739
rect 20303 48705 20312 48739
rect 20260 48696 20312 48705
rect 20996 48739 21048 48748
rect 20996 48705 21005 48739
rect 21005 48705 21039 48739
rect 21039 48705 21048 48739
rect 20996 48696 21048 48705
rect 27988 48764 28040 48816
rect 29092 48807 29144 48816
rect 29092 48773 29101 48807
rect 29101 48773 29135 48807
rect 29135 48773 29144 48807
rect 29092 48764 29144 48773
rect 20536 48628 20588 48680
rect 26516 48696 26568 48748
rect 27896 48696 27948 48748
rect 28724 48696 28776 48748
rect 29552 48764 29604 48816
rect 30288 48764 30340 48816
rect 41420 48832 41472 48884
rect 42616 48832 42668 48884
rect 43904 48875 43956 48884
rect 34796 48739 34848 48748
rect 34796 48705 34805 48739
rect 34805 48705 34839 48739
rect 34839 48705 34848 48739
rect 34796 48696 34848 48705
rect 37372 48696 37424 48748
rect 43168 48764 43220 48816
rect 43904 48841 43913 48875
rect 43913 48841 43947 48875
rect 43947 48841 43956 48875
rect 43904 48832 43956 48841
rect 45928 48875 45980 48884
rect 45928 48841 45937 48875
rect 45937 48841 45971 48875
rect 45971 48841 45980 48875
rect 45928 48832 45980 48841
rect 46020 48875 46072 48884
rect 46020 48841 46029 48875
rect 46029 48841 46063 48875
rect 46063 48841 46072 48875
rect 46940 48875 46992 48884
rect 46020 48832 46072 48841
rect 46940 48841 46949 48875
rect 46949 48841 46983 48875
rect 46983 48841 46992 48875
rect 46940 48832 46992 48841
rect 24860 48628 24912 48680
rect 27620 48628 27672 48680
rect 28448 48628 28500 48680
rect 34704 48628 34756 48680
rect 30104 48560 30156 48612
rect 14096 48492 14148 48544
rect 20444 48535 20496 48544
rect 20444 48501 20453 48535
rect 20453 48501 20487 48535
rect 20487 48501 20496 48535
rect 20444 48492 20496 48501
rect 25412 48535 25464 48544
rect 25412 48501 25421 48535
rect 25421 48501 25455 48535
rect 25455 48501 25464 48535
rect 25412 48492 25464 48501
rect 30012 48492 30064 48544
rect 33416 48492 33468 48544
rect 37556 48492 37608 48544
rect 37924 48492 37976 48544
rect 40224 48628 40276 48680
rect 41328 48671 41380 48680
rect 41328 48637 41337 48671
rect 41337 48637 41371 48671
rect 41371 48637 41380 48671
rect 41328 48628 41380 48637
rect 41604 48696 41656 48748
rect 42984 48739 43036 48748
rect 41788 48628 41840 48680
rect 42984 48705 42993 48739
rect 42993 48705 43027 48739
rect 43027 48705 43036 48739
rect 42984 48696 43036 48705
rect 43076 48671 43128 48680
rect 43076 48637 43085 48671
rect 43085 48637 43119 48671
rect 43119 48637 43128 48671
rect 43076 48628 43128 48637
rect 43720 48739 43772 48748
rect 43720 48705 43729 48739
rect 43729 48705 43763 48739
rect 43763 48705 43772 48739
rect 43720 48696 43772 48705
rect 45744 48764 45796 48816
rect 48136 48832 48188 48884
rect 51632 48875 51684 48884
rect 51632 48841 51641 48875
rect 51641 48841 51675 48875
rect 51675 48841 51684 48875
rect 51632 48832 51684 48841
rect 47584 48807 47636 48816
rect 45100 48696 45152 48748
rect 46204 48739 46256 48748
rect 46204 48705 46213 48739
rect 46213 48705 46247 48739
rect 46247 48705 46256 48739
rect 46204 48696 46256 48705
rect 47584 48773 47593 48807
rect 47593 48773 47627 48807
rect 47627 48773 47636 48807
rect 47584 48764 47636 48773
rect 47676 48764 47728 48816
rect 41420 48560 41472 48612
rect 45652 48603 45704 48612
rect 45652 48569 45661 48603
rect 45661 48569 45695 48603
rect 45695 48569 45704 48603
rect 45652 48560 45704 48569
rect 47584 48628 47636 48680
rect 50160 48696 50212 48748
rect 51356 48696 51408 48748
rect 40684 48492 40736 48544
rect 40960 48492 41012 48544
rect 45192 48492 45244 48544
rect 46204 48492 46256 48544
rect 47032 48492 47084 48544
rect 47952 48535 48004 48544
rect 47952 48501 47961 48535
rect 47961 48501 47995 48535
rect 47995 48501 48004 48535
rect 47952 48492 48004 48501
rect 49424 48492 49476 48544
rect 49700 48535 49752 48544
rect 49700 48501 49709 48535
rect 49709 48501 49743 48535
rect 49743 48501 49752 48535
rect 49700 48492 49752 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 65654 48390 65706 48442
rect 65718 48390 65770 48442
rect 65782 48390 65834 48442
rect 65846 48390 65898 48442
rect 65910 48390 65962 48442
rect 19800 48331 19852 48340
rect 19800 48297 19809 48331
rect 19809 48297 19843 48331
rect 19843 48297 19852 48331
rect 19800 48288 19852 48297
rect 19984 48331 20036 48340
rect 19984 48297 19993 48331
rect 19993 48297 20027 48331
rect 20027 48297 20036 48331
rect 19984 48288 20036 48297
rect 20444 48195 20496 48204
rect 1676 48084 1728 48136
rect 13360 48084 13412 48136
rect 14464 48127 14516 48136
rect 14464 48093 14473 48127
rect 14473 48093 14507 48127
rect 14507 48093 14516 48127
rect 14464 48084 14516 48093
rect 15292 48084 15344 48136
rect 20444 48161 20453 48195
rect 20453 48161 20487 48195
rect 20487 48161 20496 48195
rect 20444 48152 20496 48161
rect 16764 48084 16816 48136
rect 17408 48084 17460 48136
rect 20720 48127 20772 48136
rect 20720 48093 20754 48127
rect 20754 48093 20772 48127
rect 20720 48084 20772 48093
rect 17960 48016 18012 48068
rect 18052 48016 18104 48068
rect 23296 48127 23348 48136
rect 23296 48093 23305 48127
rect 23305 48093 23339 48127
rect 23339 48093 23348 48127
rect 23296 48084 23348 48093
rect 12716 47991 12768 48000
rect 12716 47957 12725 47991
rect 12725 47957 12759 47991
rect 12759 47957 12768 47991
rect 12716 47948 12768 47957
rect 14188 47948 14240 48000
rect 15016 47991 15068 48000
rect 15016 47957 15025 47991
rect 15025 47957 15059 47991
rect 15059 47957 15068 47991
rect 15016 47948 15068 47957
rect 16304 47948 16356 48000
rect 17040 47991 17092 48000
rect 17040 47957 17049 47991
rect 17049 47957 17083 47991
rect 17083 47957 17092 47991
rect 17040 47948 17092 47957
rect 20168 47948 20220 48000
rect 23664 48016 23716 48068
rect 24308 48084 24360 48136
rect 25412 48084 25464 48136
rect 29368 48220 29420 48272
rect 30288 48220 30340 48272
rect 30380 48220 30432 48272
rect 31576 48220 31628 48272
rect 32680 48220 32732 48272
rect 32864 48263 32916 48272
rect 32864 48229 32873 48263
rect 32873 48229 32907 48263
rect 32907 48229 32916 48263
rect 32864 48220 32916 48229
rect 32956 48220 33008 48272
rect 37372 48263 37424 48272
rect 37372 48229 37381 48263
rect 37381 48229 37415 48263
rect 37415 48229 37424 48263
rect 37372 48220 37424 48229
rect 41328 48288 41380 48340
rect 41880 48288 41932 48340
rect 39488 48220 39540 48272
rect 41788 48263 41840 48272
rect 41788 48229 41797 48263
rect 41797 48229 41831 48263
rect 41831 48229 41840 48263
rect 41788 48220 41840 48229
rect 23296 47948 23348 48000
rect 24860 47948 24912 48000
rect 25872 47948 25924 48000
rect 27528 48084 27580 48136
rect 33692 48195 33744 48204
rect 33692 48161 33701 48195
rect 33701 48161 33735 48195
rect 33735 48161 33744 48195
rect 33692 48152 33744 48161
rect 30564 48084 30616 48136
rect 27436 48016 27488 48068
rect 32680 48084 32732 48136
rect 33140 48127 33192 48136
rect 33140 48093 33149 48127
rect 33149 48093 33183 48127
rect 33183 48093 33192 48127
rect 33140 48084 33192 48093
rect 32496 48016 32548 48068
rect 33232 48016 33284 48068
rect 26516 47948 26568 48000
rect 27160 47991 27212 48000
rect 27160 47957 27169 47991
rect 27169 47957 27203 47991
rect 27203 47957 27212 47991
rect 27160 47948 27212 47957
rect 29184 47948 29236 48000
rect 30196 47948 30248 48000
rect 31116 47991 31168 48000
rect 31116 47957 31125 47991
rect 31125 47957 31159 47991
rect 31159 47957 31168 47991
rect 31116 47948 31168 47957
rect 32956 47948 33008 48000
rect 33968 48152 34020 48204
rect 40132 48152 40184 48204
rect 41512 48152 41564 48204
rect 41696 48152 41748 48204
rect 43168 48220 43220 48272
rect 43720 48288 43772 48340
rect 43904 48288 43956 48340
rect 46020 48288 46072 48340
rect 47032 48263 47084 48272
rect 47032 48229 47041 48263
rect 47041 48229 47075 48263
rect 47075 48229 47084 48263
rect 47032 48220 47084 48229
rect 43260 48152 43312 48204
rect 45008 48152 45060 48204
rect 34428 48084 34480 48136
rect 35624 48084 35676 48136
rect 36176 48084 36228 48136
rect 33876 48059 33928 48068
rect 33876 48025 33885 48059
rect 33885 48025 33919 48059
rect 33919 48025 33928 48059
rect 33876 48016 33928 48025
rect 37280 48084 37332 48136
rect 40040 48127 40092 48136
rect 40040 48093 40049 48127
rect 40049 48093 40083 48127
rect 40083 48093 40092 48127
rect 40040 48084 40092 48093
rect 40224 48127 40276 48136
rect 40224 48093 40233 48127
rect 40233 48093 40267 48127
rect 40267 48093 40276 48127
rect 40224 48084 40276 48093
rect 44272 48127 44324 48136
rect 37924 48016 37976 48068
rect 38016 48016 38068 48068
rect 40684 48016 40736 48068
rect 41328 48016 41380 48068
rect 41604 48059 41656 48068
rect 41604 48025 41629 48059
rect 41629 48025 41656 48059
rect 43076 48059 43128 48068
rect 41604 48016 41656 48025
rect 43076 48025 43085 48059
rect 43085 48025 43119 48059
rect 43119 48025 43128 48059
rect 43076 48016 43128 48025
rect 44272 48093 44281 48127
rect 44281 48093 44315 48127
rect 44315 48093 44324 48127
rect 44272 48084 44324 48093
rect 44456 48127 44508 48136
rect 44456 48093 44465 48127
rect 44465 48093 44499 48127
rect 44499 48093 44508 48127
rect 44456 48084 44508 48093
rect 44916 48084 44968 48136
rect 47124 48152 47176 48204
rect 45284 48127 45336 48136
rect 45284 48093 45293 48127
rect 45293 48093 45327 48127
rect 45327 48093 45336 48127
rect 45284 48084 45336 48093
rect 45468 48084 45520 48136
rect 45652 48016 45704 48068
rect 47952 48084 48004 48136
rect 48688 48084 48740 48136
rect 49148 48016 49200 48068
rect 49424 48127 49476 48136
rect 49424 48093 49433 48127
rect 49433 48093 49467 48127
rect 49467 48093 49476 48127
rect 49424 48084 49476 48093
rect 49700 48152 49752 48204
rect 67732 48059 67784 48068
rect 39856 47991 39908 48000
rect 39856 47957 39865 47991
rect 39865 47957 39899 47991
rect 39899 47957 39908 47991
rect 39856 47948 39908 47957
rect 42616 47948 42668 48000
rect 47216 47991 47268 48000
rect 47216 47957 47225 47991
rect 47225 47957 47259 47991
rect 47259 47957 47268 47991
rect 47216 47948 47268 47957
rect 47492 47948 47544 48000
rect 67732 48025 67741 48059
rect 67741 48025 67775 48059
rect 67775 48025 67784 48059
rect 67732 48016 67784 48025
rect 50160 47948 50212 48000
rect 67824 47991 67876 48000
rect 67824 47957 67833 47991
rect 67833 47957 67867 47991
rect 67867 47957 67876 47991
rect 67824 47948 67876 47957
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 17408 47787 17460 47796
rect 17408 47753 17417 47787
rect 17417 47753 17451 47787
rect 17451 47753 17460 47787
rect 17408 47744 17460 47753
rect 17960 47744 18012 47796
rect 24308 47787 24360 47796
rect 12716 47676 12768 47728
rect 15016 47676 15068 47728
rect 1676 47651 1728 47660
rect 1676 47617 1685 47651
rect 1685 47617 1719 47651
rect 1719 47617 1728 47651
rect 1676 47608 1728 47617
rect 14188 47651 14240 47660
rect 14188 47617 14197 47651
rect 14197 47617 14231 47651
rect 14231 47617 14240 47651
rect 14188 47608 14240 47617
rect 17316 47608 17368 47660
rect 18052 47651 18104 47660
rect 18052 47617 18061 47651
rect 18061 47617 18095 47651
rect 18095 47617 18104 47651
rect 18052 47608 18104 47617
rect 24308 47753 24317 47787
rect 24317 47753 24351 47787
rect 24351 47753 24360 47787
rect 24308 47744 24360 47753
rect 27528 47787 27580 47796
rect 27528 47753 27537 47787
rect 27537 47753 27571 47787
rect 27571 47753 27580 47787
rect 27528 47744 27580 47753
rect 2412 47540 2464 47592
rect 2780 47583 2832 47592
rect 2780 47549 2789 47583
rect 2789 47549 2823 47583
rect 2823 47549 2832 47583
rect 2780 47540 2832 47549
rect 12164 47583 12216 47592
rect 12164 47549 12173 47583
rect 12173 47549 12207 47583
rect 12207 47549 12216 47583
rect 12164 47540 12216 47549
rect 17684 47540 17736 47592
rect 15568 47515 15620 47524
rect 15568 47481 15577 47515
rect 15577 47481 15611 47515
rect 15611 47481 15620 47515
rect 18880 47583 18932 47592
rect 18880 47549 18914 47583
rect 18914 47549 18932 47583
rect 18880 47540 18932 47549
rect 19064 47583 19116 47592
rect 19064 47549 19073 47583
rect 19073 47549 19107 47583
rect 19107 47549 19116 47583
rect 19064 47540 19116 47549
rect 20996 47540 21048 47592
rect 25872 47676 25924 47728
rect 23112 47608 23164 47660
rect 24308 47651 24360 47660
rect 24308 47617 24317 47651
rect 24317 47617 24351 47651
rect 24351 47617 24360 47651
rect 24308 47608 24360 47617
rect 26240 47651 26292 47660
rect 26240 47617 26249 47651
rect 26249 47617 26283 47651
rect 26283 47617 26292 47651
rect 27804 47676 27856 47728
rect 26240 47608 26292 47617
rect 27436 47608 27488 47660
rect 33784 47744 33836 47796
rect 33968 47744 34020 47796
rect 35440 47744 35492 47796
rect 35808 47787 35860 47796
rect 35808 47753 35817 47787
rect 35817 47753 35851 47787
rect 35851 47753 35860 47787
rect 35808 47744 35860 47753
rect 35992 47744 36044 47796
rect 67824 47744 67876 47796
rect 28540 47719 28592 47728
rect 28540 47685 28549 47719
rect 28549 47685 28583 47719
rect 28583 47685 28592 47719
rect 28540 47676 28592 47685
rect 29092 47676 29144 47728
rect 28448 47651 28500 47660
rect 25872 47540 25924 47592
rect 28448 47617 28457 47651
rect 28457 47617 28491 47651
rect 28491 47617 28500 47651
rect 28448 47608 28500 47617
rect 28908 47540 28960 47592
rect 31116 47676 31168 47728
rect 30196 47651 30248 47660
rect 30196 47617 30205 47651
rect 30205 47617 30239 47651
rect 30239 47617 30248 47651
rect 30196 47608 30248 47617
rect 34704 47676 34756 47728
rect 32864 47651 32916 47660
rect 32864 47617 32898 47651
rect 32898 47617 32916 47651
rect 32864 47608 32916 47617
rect 33140 47608 33192 47660
rect 33784 47608 33836 47660
rect 35532 47676 35584 47728
rect 36360 47676 36412 47728
rect 35624 47608 35676 47660
rect 37832 47651 37884 47660
rect 15568 47472 15620 47481
rect 18236 47472 18288 47524
rect 33692 47540 33744 47592
rect 34336 47540 34388 47592
rect 35624 47472 35676 47524
rect 13544 47447 13596 47456
rect 13544 47413 13553 47447
rect 13553 47413 13587 47447
rect 13587 47413 13596 47447
rect 13544 47404 13596 47413
rect 18880 47404 18932 47456
rect 21088 47404 21140 47456
rect 23664 47447 23716 47456
rect 23664 47413 23673 47447
rect 23673 47413 23707 47447
rect 23707 47413 23716 47447
rect 23664 47404 23716 47413
rect 24768 47404 24820 47456
rect 26424 47404 26476 47456
rect 29460 47447 29512 47456
rect 29460 47413 29469 47447
rect 29469 47413 29503 47447
rect 29503 47413 29512 47447
rect 29460 47404 29512 47413
rect 30196 47404 30248 47456
rect 33600 47404 33652 47456
rect 34612 47447 34664 47456
rect 34612 47413 34621 47447
rect 34621 47413 34655 47447
rect 34655 47413 34664 47447
rect 34612 47404 34664 47413
rect 34796 47404 34848 47456
rect 35440 47404 35492 47456
rect 37832 47617 37841 47651
rect 37841 47617 37875 47651
rect 37875 47617 37884 47651
rect 37832 47608 37884 47617
rect 38752 47404 38804 47456
rect 39396 47651 39448 47660
rect 39396 47617 39405 47651
rect 39405 47617 39439 47651
rect 39439 47617 39448 47651
rect 39396 47608 39448 47617
rect 39948 47608 40000 47660
rect 40960 47651 41012 47660
rect 39672 47540 39724 47592
rect 40960 47617 40969 47651
rect 40969 47617 41003 47651
rect 41003 47617 41012 47651
rect 40960 47608 41012 47617
rect 42616 47676 42668 47728
rect 43260 47719 43312 47728
rect 43260 47685 43269 47719
rect 43269 47685 43303 47719
rect 43303 47685 43312 47719
rect 43260 47676 43312 47685
rect 47952 47676 48004 47728
rect 48688 47719 48740 47728
rect 48688 47685 48697 47719
rect 48697 47685 48731 47719
rect 48731 47685 48740 47719
rect 48688 47676 48740 47685
rect 49148 47676 49200 47728
rect 49700 47676 49752 47728
rect 50160 47676 50212 47728
rect 41420 47651 41472 47660
rect 41420 47617 41429 47651
rect 41429 47617 41463 47651
rect 41463 47617 41472 47651
rect 41420 47608 41472 47617
rect 44916 47651 44968 47660
rect 40960 47472 41012 47524
rect 43076 47540 43128 47592
rect 43628 47583 43680 47592
rect 43628 47549 43637 47583
rect 43637 47549 43671 47583
rect 43671 47549 43680 47583
rect 43628 47540 43680 47549
rect 41328 47472 41380 47524
rect 44916 47617 44925 47651
rect 44925 47617 44959 47651
rect 44959 47617 44968 47651
rect 44916 47608 44968 47617
rect 45652 47608 45704 47660
rect 48596 47608 48648 47660
rect 50620 47651 50672 47660
rect 44272 47540 44324 47592
rect 46296 47540 46348 47592
rect 49792 47540 49844 47592
rect 50620 47617 50629 47651
rect 50629 47617 50663 47651
rect 50663 47617 50672 47651
rect 50620 47608 50672 47617
rect 51448 47608 51500 47660
rect 51632 47651 51684 47660
rect 51632 47617 51641 47651
rect 51641 47617 51675 47651
rect 51675 47617 51684 47651
rect 51632 47608 51684 47617
rect 50804 47540 50856 47592
rect 40040 47404 40092 47456
rect 40684 47447 40736 47456
rect 40684 47413 40693 47447
rect 40693 47413 40727 47447
rect 40727 47413 40736 47447
rect 40684 47404 40736 47413
rect 41788 47404 41840 47456
rect 43168 47404 43220 47456
rect 44640 47472 44692 47524
rect 44364 47404 44416 47456
rect 45192 47447 45244 47456
rect 45192 47413 45201 47447
rect 45201 47413 45235 47447
rect 45235 47413 45244 47447
rect 45192 47404 45244 47413
rect 51724 47404 51776 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 65654 47302 65706 47354
rect 65718 47302 65770 47354
rect 65782 47302 65834 47354
rect 65846 47302 65898 47354
rect 65910 47302 65962 47354
rect 2412 47243 2464 47252
rect 2412 47209 2421 47243
rect 2421 47209 2455 47243
rect 2455 47209 2464 47243
rect 2412 47200 2464 47209
rect 12164 47200 12216 47252
rect 13360 47243 13412 47252
rect 13360 47209 13369 47243
rect 13369 47209 13403 47243
rect 13403 47209 13412 47243
rect 13360 47200 13412 47209
rect 15292 47243 15344 47252
rect 15292 47209 15301 47243
rect 15301 47209 15335 47243
rect 15335 47209 15344 47243
rect 15292 47200 15344 47209
rect 17684 47243 17736 47252
rect 17684 47209 17693 47243
rect 17693 47209 17727 47243
rect 17727 47209 17736 47243
rect 17684 47200 17736 47209
rect 23112 47243 23164 47252
rect 23112 47209 23121 47243
rect 23121 47209 23155 47243
rect 23155 47209 23164 47243
rect 23112 47200 23164 47209
rect 27804 47243 27856 47252
rect 27804 47209 27813 47243
rect 27813 47209 27847 47243
rect 27847 47209 27856 47243
rect 27804 47200 27856 47209
rect 30380 47243 30432 47252
rect 30380 47209 30389 47243
rect 30389 47209 30423 47243
rect 30423 47209 30432 47243
rect 30380 47200 30432 47209
rect 30564 47243 30616 47252
rect 30564 47209 30573 47243
rect 30573 47209 30607 47243
rect 30607 47209 30616 47243
rect 30564 47200 30616 47209
rect 32956 47200 33008 47252
rect 33968 47243 34020 47252
rect 33968 47209 33977 47243
rect 33977 47209 34011 47243
rect 34011 47209 34020 47243
rect 33968 47200 34020 47209
rect 14096 47132 14148 47184
rect 30288 47132 30340 47184
rect 38016 47200 38068 47252
rect 39396 47200 39448 47252
rect 40224 47243 40276 47252
rect 34796 47132 34848 47184
rect 13544 47064 13596 47116
rect 15568 47064 15620 47116
rect 16304 47107 16356 47116
rect 16304 47073 16313 47107
rect 16313 47073 16347 47107
rect 16347 47073 16356 47107
rect 16304 47064 16356 47073
rect 20168 47064 20220 47116
rect 26424 47107 26476 47116
rect 26424 47073 26433 47107
rect 26433 47073 26467 47107
rect 26467 47073 26476 47107
rect 26424 47064 26476 47073
rect 29276 47064 29328 47116
rect 33600 47064 33652 47116
rect 34336 47064 34388 47116
rect 37832 47132 37884 47184
rect 35440 47064 35492 47116
rect 2320 47039 2372 47048
rect 2320 47005 2329 47039
rect 2329 47005 2363 47039
rect 2363 47005 2372 47039
rect 2320 46996 2372 47005
rect 6828 46996 6880 47048
rect 12624 46996 12676 47048
rect 13268 46996 13320 47048
rect 15292 46996 15344 47048
rect 17040 46996 17092 47048
rect 20812 46996 20864 47048
rect 20996 47039 21048 47048
rect 20996 47005 21005 47039
rect 21005 47005 21039 47039
rect 21039 47005 21048 47039
rect 20996 46996 21048 47005
rect 21824 47039 21876 47048
rect 21824 47005 21833 47039
rect 21833 47005 21867 47039
rect 21867 47005 21876 47039
rect 21824 46996 21876 47005
rect 23296 47039 23348 47048
rect 23296 47005 23305 47039
rect 23305 47005 23339 47039
rect 23339 47005 23348 47039
rect 23296 46996 23348 47005
rect 27160 46996 27212 47048
rect 31576 46996 31628 47048
rect 32496 47039 32548 47048
rect 32496 47005 32505 47039
rect 32505 47005 32539 47039
rect 32539 47005 32548 47039
rect 32496 46996 32548 47005
rect 35808 47064 35860 47116
rect 25596 46928 25648 46980
rect 30196 46971 30248 46980
rect 30196 46937 30205 46971
rect 30205 46937 30239 46971
rect 30239 46937 30248 46971
rect 30196 46928 30248 46937
rect 30288 46928 30340 46980
rect 30564 46928 30616 46980
rect 33508 46928 33560 46980
rect 33784 46971 33836 46980
rect 33784 46937 33793 46971
rect 33793 46937 33827 46971
rect 33827 46937 33836 46971
rect 33784 46928 33836 46937
rect 35532 46928 35584 46980
rect 36452 47039 36504 47048
rect 36452 47005 36461 47039
rect 36461 47005 36495 47039
rect 36495 47005 36504 47039
rect 36452 46996 36504 47005
rect 36728 47039 36780 47048
rect 36728 47005 36737 47039
rect 36737 47005 36771 47039
rect 36771 47005 36780 47039
rect 36728 46996 36780 47005
rect 36360 46928 36412 46980
rect 37280 46928 37332 46980
rect 19984 46860 20036 46912
rect 20812 46903 20864 46912
rect 20812 46869 20821 46903
rect 20821 46869 20855 46903
rect 20855 46869 20864 46903
rect 20812 46860 20864 46869
rect 24032 46860 24084 46912
rect 24860 46860 24912 46912
rect 28908 46903 28960 46912
rect 28908 46869 28917 46903
rect 28917 46869 28951 46903
rect 28951 46869 28960 46903
rect 28908 46860 28960 46869
rect 31852 46903 31904 46912
rect 31852 46869 31861 46903
rect 31861 46869 31895 46903
rect 31895 46869 31904 46903
rect 31852 46860 31904 46869
rect 32036 46860 32088 46912
rect 38016 47039 38068 47048
rect 38016 47005 38025 47039
rect 38025 47005 38059 47039
rect 38059 47005 38068 47039
rect 38016 46996 38068 47005
rect 38108 46996 38160 47048
rect 38936 47039 38988 47048
rect 38936 47005 38945 47039
rect 38945 47005 38979 47039
rect 38979 47005 38988 47039
rect 38936 46996 38988 47005
rect 40224 47209 40233 47243
rect 40233 47209 40267 47243
rect 40267 47209 40276 47243
rect 40224 47200 40276 47209
rect 44364 47200 44416 47252
rect 46112 47200 46164 47252
rect 46296 47243 46348 47252
rect 46296 47209 46305 47243
rect 46305 47209 46339 47243
rect 46339 47209 46348 47243
rect 46296 47200 46348 47209
rect 46664 47243 46716 47252
rect 46664 47209 46673 47243
rect 46673 47209 46707 47243
rect 46707 47209 46716 47243
rect 46664 47200 46716 47209
rect 51448 47200 51500 47252
rect 41696 47132 41748 47184
rect 40132 47064 40184 47116
rect 40960 47064 41012 47116
rect 45836 47064 45888 47116
rect 66996 47064 67048 47116
rect 67180 47064 67232 47116
rect 44456 46996 44508 47048
rect 44916 46996 44968 47048
rect 45652 47039 45704 47048
rect 37924 46928 37976 46980
rect 39948 46928 40000 46980
rect 40040 46971 40092 46980
rect 40040 46937 40065 46971
rect 40065 46937 40092 46971
rect 40040 46928 40092 46937
rect 43444 46928 43496 46980
rect 45652 47005 45661 47039
rect 45661 47005 45695 47039
rect 45695 47005 45704 47039
rect 45652 46996 45704 47005
rect 46388 47039 46440 47048
rect 46388 47005 46397 47039
rect 46397 47005 46431 47039
rect 46431 47005 46440 47039
rect 46388 46996 46440 47005
rect 51724 46996 51776 47048
rect 66260 46996 66312 47048
rect 51356 46928 51408 46980
rect 58716 46928 58768 46980
rect 67088 46928 67140 46980
rect 46388 46860 46440 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 22100 46656 22152 46708
rect 17316 46588 17368 46640
rect 20812 46588 20864 46640
rect 28632 46656 28684 46708
rect 32956 46656 33008 46708
rect 35624 46656 35676 46708
rect 36268 46656 36320 46708
rect 42616 46699 42668 46708
rect 42616 46665 42625 46699
rect 42625 46665 42659 46699
rect 42659 46665 42668 46699
rect 42616 46656 42668 46665
rect 43168 46699 43220 46708
rect 43168 46665 43177 46699
rect 43177 46665 43211 46699
rect 43211 46665 43220 46699
rect 43168 46656 43220 46665
rect 45560 46656 45612 46708
rect 47584 46656 47636 46708
rect 50804 46699 50856 46708
rect 50804 46665 50813 46699
rect 50813 46665 50847 46699
rect 50847 46665 50856 46699
rect 50804 46656 50856 46665
rect 51632 46656 51684 46708
rect 1860 46563 1912 46572
rect 1860 46529 1869 46563
rect 1869 46529 1903 46563
rect 1903 46529 1912 46563
rect 1860 46520 1912 46529
rect 17408 46563 17460 46572
rect 17408 46529 17417 46563
rect 17417 46529 17451 46563
rect 17451 46529 17460 46563
rect 17408 46520 17460 46529
rect 17500 46563 17552 46572
rect 17500 46529 17509 46563
rect 17509 46529 17543 46563
rect 17543 46529 17552 46563
rect 17500 46520 17552 46529
rect 18972 46520 19024 46572
rect 19984 46520 20036 46572
rect 20904 46520 20956 46572
rect 22284 46520 22336 46572
rect 24032 46563 24084 46572
rect 24032 46529 24041 46563
rect 24041 46529 24075 46563
rect 24075 46529 24084 46563
rect 24032 46520 24084 46529
rect 24952 46563 25004 46572
rect 24952 46529 24961 46563
rect 24961 46529 24995 46563
rect 24995 46529 25004 46563
rect 24952 46520 25004 46529
rect 27988 46520 28040 46572
rect 28908 46520 28960 46572
rect 29276 46563 29328 46572
rect 29276 46529 29285 46563
rect 29285 46529 29319 46563
rect 29319 46529 29328 46563
rect 29276 46520 29328 46529
rect 30012 46563 30064 46572
rect 30012 46529 30021 46563
rect 30021 46529 30055 46563
rect 30055 46529 30064 46563
rect 30012 46520 30064 46529
rect 30932 46563 30984 46572
rect 30932 46529 30941 46563
rect 30941 46529 30975 46563
rect 30975 46529 30984 46563
rect 30932 46520 30984 46529
rect 24768 46452 24820 46504
rect 25044 46495 25096 46504
rect 25044 46461 25078 46495
rect 25078 46461 25096 46495
rect 25044 46452 25096 46461
rect 26056 46452 26108 46504
rect 33416 46520 33468 46572
rect 35900 46520 35952 46572
rect 36728 46520 36780 46572
rect 37280 46520 37332 46572
rect 38568 46563 38620 46572
rect 38568 46529 38577 46563
rect 38577 46529 38611 46563
rect 38611 46529 38620 46563
rect 38568 46520 38620 46529
rect 40224 46588 40276 46640
rect 40684 46520 40736 46572
rect 41696 46563 41748 46572
rect 41696 46529 41705 46563
rect 41705 46529 41739 46563
rect 41739 46529 41748 46563
rect 41696 46520 41748 46529
rect 42064 46588 42116 46640
rect 47124 46588 47176 46640
rect 47216 46588 47268 46640
rect 48044 46588 48096 46640
rect 49700 46631 49752 46640
rect 49700 46597 49734 46631
rect 49734 46597 49752 46631
rect 49700 46588 49752 46597
rect 42432 46520 42484 46572
rect 43904 46520 43956 46572
rect 44364 46520 44416 46572
rect 45652 46563 45704 46572
rect 31852 46452 31904 46504
rect 32496 46452 32548 46504
rect 32772 46495 32824 46504
rect 32772 46461 32781 46495
rect 32781 46461 32815 46495
rect 32815 46461 32824 46495
rect 32772 46452 32824 46461
rect 32864 46452 32916 46504
rect 35348 46452 35400 46504
rect 38200 46452 38252 46504
rect 39948 46452 40000 46504
rect 2044 46427 2096 46436
rect 2044 46393 2053 46427
rect 2053 46393 2087 46427
rect 2087 46393 2096 46427
rect 2044 46384 2096 46393
rect 18512 46316 18564 46368
rect 19248 46359 19300 46368
rect 19248 46325 19257 46359
rect 19257 46325 19291 46359
rect 19291 46325 19300 46359
rect 19248 46316 19300 46325
rect 19708 46316 19760 46368
rect 21640 46316 21692 46368
rect 21916 46316 21968 46368
rect 25688 46316 25740 46368
rect 26332 46384 26384 46436
rect 33784 46384 33836 46436
rect 38292 46384 38344 46436
rect 39028 46384 39080 46436
rect 43444 46427 43496 46436
rect 43444 46393 43453 46427
rect 43453 46393 43487 46427
rect 43487 46393 43496 46427
rect 43444 46384 43496 46393
rect 43536 46427 43588 46436
rect 43536 46393 43545 46427
rect 43545 46393 43579 46427
rect 43579 46393 43588 46427
rect 43536 46384 43588 46393
rect 28632 46359 28684 46368
rect 28632 46325 28641 46359
rect 28641 46325 28675 46359
rect 28675 46325 28684 46359
rect 28632 46316 28684 46325
rect 29000 46316 29052 46368
rect 29368 46316 29420 46368
rect 29920 46316 29972 46368
rect 30748 46359 30800 46368
rect 30748 46325 30757 46359
rect 30757 46325 30791 46359
rect 30791 46325 30800 46359
rect 30748 46316 30800 46325
rect 38660 46316 38712 46368
rect 39120 46316 39172 46368
rect 40132 46316 40184 46368
rect 42156 46316 42208 46368
rect 45652 46529 45661 46563
rect 45661 46529 45695 46563
rect 45695 46529 45704 46563
rect 45652 46520 45704 46529
rect 51448 46520 51500 46572
rect 51724 46563 51776 46572
rect 51724 46529 51733 46563
rect 51733 46529 51767 46563
rect 51767 46529 51776 46563
rect 51724 46520 51776 46529
rect 66260 46588 66312 46640
rect 45836 46452 45888 46504
rect 49424 46495 49476 46504
rect 49424 46461 49433 46495
rect 49433 46461 49467 46495
rect 49467 46461 49476 46495
rect 49424 46452 49476 46461
rect 67364 46452 67416 46504
rect 67548 46495 67600 46504
rect 67548 46461 67557 46495
rect 67557 46461 67591 46495
rect 67591 46461 67600 46495
rect 67548 46452 67600 46461
rect 45100 46316 45152 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 65654 46214 65706 46266
rect 65718 46214 65770 46266
rect 65782 46214 65834 46266
rect 65846 46214 65898 46266
rect 65910 46214 65962 46266
rect 17408 46112 17460 46164
rect 19984 46112 20036 46164
rect 20996 46044 21048 46096
rect 19248 45976 19300 46028
rect 24032 46112 24084 46164
rect 25688 46112 25740 46164
rect 26056 46112 26108 46164
rect 33508 46112 33560 46164
rect 36176 46112 36228 46164
rect 42432 46112 42484 46164
rect 43444 46155 43496 46164
rect 43444 46121 43453 46155
rect 43453 46121 43487 46155
rect 43487 46121 43496 46155
rect 43444 46112 43496 46121
rect 45284 46112 45336 46164
rect 45652 46112 45704 46164
rect 49424 46112 49476 46164
rect 66812 46112 66864 46164
rect 67180 46112 67232 46164
rect 67364 46155 67416 46164
rect 67364 46121 67373 46155
rect 67373 46121 67407 46155
rect 67407 46121 67416 46155
rect 67364 46112 67416 46121
rect 45100 46087 45152 46096
rect 45100 46053 45109 46087
rect 45109 46053 45143 46087
rect 45143 46053 45152 46087
rect 45100 46044 45152 46053
rect 21640 46019 21692 46028
rect 21640 45985 21649 46019
rect 21649 45985 21683 46019
rect 21683 45985 21692 46019
rect 21640 45976 21692 45985
rect 13544 45908 13596 45960
rect 14464 45951 14516 45960
rect 14464 45917 14473 45951
rect 14473 45917 14507 45951
rect 14507 45917 14516 45951
rect 14464 45908 14516 45917
rect 15476 45908 15528 45960
rect 16580 45908 16632 45960
rect 18512 45951 18564 45960
rect 18512 45917 18521 45951
rect 18521 45917 18555 45951
rect 18555 45917 18564 45951
rect 18512 45908 18564 45917
rect 18972 45908 19024 45960
rect 21916 45951 21968 45960
rect 12992 45815 13044 45824
rect 12992 45781 13001 45815
rect 13001 45781 13035 45815
rect 13035 45781 13044 45815
rect 12992 45772 13044 45781
rect 14648 45815 14700 45824
rect 14648 45781 14657 45815
rect 14657 45781 14691 45815
rect 14691 45781 14700 45815
rect 14648 45772 14700 45781
rect 15200 45815 15252 45824
rect 15200 45781 15209 45815
rect 15209 45781 15243 45815
rect 15243 45781 15252 45815
rect 15200 45772 15252 45781
rect 19248 45840 19300 45892
rect 19708 45883 19760 45892
rect 19708 45849 19717 45883
rect 19717 45849 19751 45883
rect 19751 45849 19760 45883
rect 19708 45840 19760 45849
rect 20168 45840 20220 45892
rect 20536 45883 20588 45892
rect 20536 45849 20545 45883
rect 20545 45849 20579 45883
rect 20579 45849 20588 45883
rect 20536 45840 20588 45849
rect 21916 45917 21950 45951
rect 21950 45917 21968 45951
rect 21916 45908 21968 45917
rect 29920 46019 29972 46028
rect 24952 45908 25004 45960
rect 20628 45772 20680 45824
rect 20904 45815 20956 45824
rect 20904 45781 20913 45815
rect 20913 45781 20947 45815
rect 20947 45781 20956 45815
rect 20904 45772 20956 45781
rect 21640 45772 21692 45824
rect 23664 45815 23716 45824
rect 23664 45781 23673 45815
rect 23673 45781 23707 45815
rect 23707 45781 23716 45815
rect 23664 45772 23716 45781
rect 24676 45840 24728 45892
rect 25044 45840 25096 45892
rect 25780 45951 25832 45960
rect 25780 45917 25789 45951
rect 25789 45917 25823 45951
rect 25823 45917 25832 45951
rect 25780 45908 25832 45917
rect 29920 45985 29929 46019
rect 29929 45985 29963 46019
rect 29963 45985 29972 46019
rect 29920 45976 29972 45985
rect 32036 46019 32088 46028
rect 32036 45985 32045 46019
rect 32045 45985 32079 46019
rect 32079 45985 32088 46019
rect 32036 45976 32088 45985
rect 50620 46019 50672 46028
rect 25504 45840 25556 45892
rect 29828 45908 29880 45960
rect 30748 45908 30800 45960
rect 34060 45951 34112 45960
rect 28908 45840 28960 45892
rect 29368 45840 29420 45892
rect 34060 45917 34069 45951
rect 34069 45917 34103 45951
rect 34103 45917 34112 45951
rect 34060 45908 34112 45917
rect 34796 45908 34848 45960
rect 35532 45908 35584 45960
rect 25596 45772 25648 45824
rect 28356 45815 28408 45824
rect 28356 45781 28365 45815
rect 28365 45781 28399 45815
rect 28399 45781 28408 45815
rect 28356 45772 28408 45781
rect 30472 45772 30524 45824
rect 32680 45772 32732 45824
rect 34612 45840 34664 45892
rect 35624 45772 35676 45824
rect 50620 45985 50629 46019
rect 50629 45985 50663 46019
rect 50663 45985 50672 46019
rect 50620 45976 50672 45985
rect 40040 45951 40092 45960
rect 40040 45917 40049 45951
rect 40049 45917 40083 45951
rect 40083 45917 40092 45951
rect 40040 45908 40092 45917
rect 40132 45908 40184 45960
rect 42064 45951 42116 45960
rect 42064 45917 42073 45951
rect 42073 45917 42107 45951
rect 42107 45917 42116 45951
rect 42064 45908 42116 45917
rect 42156 45908 42208 45960
rect 36452 45840 36504 45892
rect 46388 45908 46440 45960
rect 48044 45951 48096 45960
rect 48044 45917 48053 45951
rect 48053 45917 48087 45951
rect 48087 45917 48096 45951
rect 48044 45908 48096 45917
rect 45836 45840 45888 45892
rect 66812 45908 66864 45960
rect 51724 45840 51776 45892
rect 37740 45772 37792 45824
rect 51448 45815 51500 45824
rect 51448 45781 51457 45815
rect 51457 45781 51491 45815
rect 51491 45781 51500 45815
rect 51448 45772 51500 45781
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 16580 45568 16632 45620
rect 12992 45500 13044 45552
rect 15200 45500 15252 45552
rect 1860 45475 1912 45484
rect 1860 45441 1869 45475
rect 1869 45441 1903 45475
rect 1903 45441 1912 45475
rect 1860 45432 1912 45441
rect 14648 45432 14700 45484
rect 16948 45432 17000 45484
rect 17408 45432 17460 45484
rect 19248 45568 19300 45620
rect 20628 45568 20680 45620
rect 22284 45611 22336 45620
rect 21364 45500 21416 45552
rect 22284 45577 22293 45611
rect 22293 45577 22327 45611
rect 22327 45577 22336 45611
rect 22284 45568 22336 45577
rect 24676 45611 24728 45620
rect 24676 45577 24685 45611
rect 24685 45577 24719 45611
rect 24719 45577 24728 45611
rect 24676 45568 24728 45577
rect 24768 45568 24820 45620
rect 29368 45568 29420 45620
rect 29828 45611 29880 45620
rect 29828 45577 29837 45611
rect 29837 45577 29871 45611
rect 29871 45577 29880 45611
rect 29828 45568 29880 45577
rect 30932 45568 30984 45620
rect 42064 45568 42116 45620
rect 18420 45475 18472 45484
rect 18420 45441 18429 45475
rect 18429 45441 18463 45475
rect 18463 45441 18472 45475
rect 18420 45432 18472 45441
rect 20076 45475 20128 45484
rect 20076 45441 20110 45475
rect 20110 45441 20128 45475
rect 20076 45432 20128 45441
rect 21272 45432 21324 45484
rect 21640 45432 21692 45484
rect 23664 45500 23716 45552
rect 24860 45500 24912 45552
rect 25596 45543 25648 45552
rect 25596 45509 25605 45543
rect 25605 45509 25639 45543
rect 25639 45509 25648 45543
rect 25596 45500 25648 45509
rect 25688 45500 25740 45552
rect 28356 45500 28408 45552
rect 28816 45500 28868 45552
rect 26976 45475 27028 45484
rect 26976 45441 26985 45475
rect 26985 45441 27019 45475
rect 27019 45441 27028 45475
rect 26976 45432 27028 45441
rect 30472 45500 30524 45552
rect 30564 45543 30616 45552
rect 30564 45509 30605 45543
rect 30605 45509 30616 45543
rect 32680 45543 32732 45552
rect 30564 45500 30616 45509
rect 32680 45509 32689 45543
rect 32689 45509 32723 45543
rect 32723 45509 32732 45543
rect 32680 45500 32732 45509
rect 34520 45500 34572 45552
rect 34704 45500 34756 45552
rect 12532 45407 12584 45416
rect 12532 45373 12541 45407
rect 12541 45373 12575 45407
rect 12575 45373 12584 45407
rect 12532 45364 12584 45373
rect 19064 45364 19116 45416
rect 19432 45364 19484 45416
rect 23296 45407 23348 45416
rect 23296 45373 23305 45407
rect 23305 45373 23339 45407
rect 23339 45373 23348 45407
rect 23296 45364 23348 45373
rect 25780 45364 25832 45416
rect 1952 45271 2004 45280
rect 1952 45237 1961 45271
rect 1961 45237 1995 45271
rect 1995 45237 2004 45271
rect 1952 45228 2004 45237
rect 13176 45228 13228 45280
rect 18236 45296 18288 45348
rect 27620 45407 27672 45416
rect 27620 45373 27629 45407
rect 27629 45373 27663 45407
rect 27663 45373 27672 45407
rect 27620 45364 27672 45373
rect 15936 45271 15988 45280
rect 15936 45237 15945 45271
rect 15945 45237 15979 45271
rect 15979 45237 15988 45271
rect 15936 45228 15988 45237
rect 18420 45228 18472 45280
rect 20536 45228 20588 45280
rect 25964 45271 26016 45280
rect 25964 45237 25973 45271
rect 25973 45237 26007 45271
rect 26007 45237 26016 45271
rect 25964 45228 26016 45237
rect 28816 45228 28868 45280
rect 35624 45475 35676 45484
rect 34060 45296 34112 45348
rect 35624 45441 35633 45475
rect 35633 45441 35667 45475
rect 35667 45441 35676 45475
rect 35624 45432 35676 45441
rect 34428 45407 34480 45416
rect 34428 45373 34437 45407
rect 34437 45373 34471 45407
rect 34471 45373 34480 45407
rect 34428 45364 34480 45373
rect 34796 45364 34848 45416
rect 37464 45500 37516 45552
rect 39856 45500 39908 45552
rect 43628 45500 43680 45552
rect 51448 45500 51500 45552
rect 37556 45475 37608 45484
rect 37556 45441 37590 45475
rect 37590 45441 37608 45475
rect 37556 45432 37608 45441
rect 41420 45432 41472 45484
rect 44916 45475 44968 45484
rect 44916 45441 44925 45475
rect 44925 45441 44959 45475
rect 44959 45441 44968 45475
rect 44916 45432 44968 45441
rect 45652 45432 45704 45484
rect 35716 45296 35768 45348
rect 32864 45271 32916 45280
rect 32864 45237 32873 45271
rect 32873 45237 32907 45271
rect 32907 45237 32916 45271
rect 32864 45228 32916 45237
rect 35440 45271 35492 45280
rect 35440 45237 35449 45271
rect 35449 45237 35483 45271
rect 35483 45237 35492 45271
rect 35440 45228 35492 45237
rect 36268 45271 36320 45280
rect 36268 45237 36277 45271
rect 36277 45237 36311 45271
rect 36311 45237 36320 45271
rect 36268 45228 36320 45237
rect 37464 45228 37516 45280
rect 38016 45228 38068 45280
rect 45744 45364 45796 45416
rect 47952 45432 48004 45484
rect 48044 45364 48096 45416
rect 50160 45407 50212 45416
rect 50160 45373 50169 45407
rect 50169 45373 50203 45407
rect 50203 45373 50212 45407
rect 50160 45364 50212 45373
rect 41512 45296 41564 45348
rect 48504 45296 48556 45348
rect 45560 45228 45612 45280
rect 47584 45271 47636 45280
rect 47584 45237 47593 45271
rect 47593 45237 47627 45271
rect 47627 45237 47636 45271
rect 47584 45228 47636 45237
rect 48320 45271 48372 45280
rect 48320 45237 48329 45271
rect 48329 45237 48363 45271
rect 48363 45237 48372 45271
rect 48320 45228 48372 45237
rect 50804 45228 50856 45280
rect 66260 45228 66312 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 65654 45126 65706 45178
rect 65718 45126 65770 45178
rect 65782 45126 65834 45178
rect 65846 45126 65898 45178
rect 65910 45126 65962 45178
rect 1952 45024 2004 45076
rect 12532 45024 12584 45076
rect 13544 45067 13596 45076
rect 13544 45033 13553 45067
rect 13553 45033 13587 45067
rect 13587 45033 13596 45067
rect 13544 45024 13596 45033
rect 15476 45067 15528 45076
rect 15476 45033 15485 45067
rect 15485 45033 15519 45067
rect 15519 45033 15528 45067
rect 15476 45024 15528 45033
rect 19432 45067 19484 45076
rect 19432 45033 19441 45067
rect 19441 45033 19475 45067
rect 19475 45033 19484 45067
rect 19432 45024 19484 45033
rect 20076 45024 20128 45076
rect 21456 45067 21508 45076
rect 21456 45033 21465 45067
rect 21465 45033 21499 45067
rect 21499 45033 21508 45067
rect 21456 45024 21508 45033
rect 25504 45024 25556 45076
rect 27620 45067 27672 45076
rect 27620 45033 27629 45067
rect 27629 45033 27663 45067
rect 27663 45033 27672 45067
rect 27620 45024 27672 45033
rect 28908 45067 28960 45076
rect 28908 45033 28917 45067
rect 28917 45033 28951 45067
rect 28951 45033 28960 45067
rect 28908 45024 28960 45033
rect 30656 45024 30708 45076
rect 37556 45024 37608 45076
rect 40040 45024 40092 45076
rect 45560 45024 45612 45076
rect 46664 45024 46716 45076
rect 50160 45067 50212 45076
rect 50160 45033 50169 45067
rect 50169 45033 50203 45067
rect 50203 45033 50212 45067
rect 50160 45024 50212 45033
rect 19892 44956 19944 45008
rect 30564 44956 30616 45008
rect 46296 44956 46348 45008
rect 13176 44931 13228 44940
rect 13176 44897 13185 44931
rect 13185 44897 13219 44931
rect 13219 44897 13228 44931
rect 13176 44888 13228 44897
rect 15936 44888 15988 44940
rect 12624 44863 12676 44872
rect 12624 44829 12633 44863
rect 12633 44829 12667 44863
rect 12667 44829 12676 44863
rect 12624 44820 12676 44829
rect 13360 44863 13412 44872
rect 13360 44829 13369 44863
rect 13369 44829 13403 44863
rect 13403 44829 13412 44863
rect 13360 44820 13412 44829
rect 15292 44863 15344 44872
rect 15292 44829 15301 44863
rect 15301 44829 15335 44863
rect 15335 44829 15344 44863
rect 15292 44820 15344 44829
rect 15568 44820 15620 44872
rect 20812 44888 20864 44940
rect 21088 44888 21140 44940
rect 20904 44820 20956 44872
rect 21824 44820 21876 44872
rect 26976 44888 27028 44940
rect 23572 44820 23624 44872
rect 25964 44863 26016 44872
rect 25964 44829 25973 44863
rect 25973 44829 26007 44863
rect 26007 44829 26016 44863
rect 25964 44820 26016 44829
rect 30012 44888 30064 44940
rect 34704 44888 34756 44940
rect 38016 44888 38068 44940
rect 28356 44820 28408 44872
rect 31116 44863 31168 44872
rect 31116 44829 31125 44863
rect 31125 44829 31159 44863
rect 31159 44829 31168 44863
rect 31116 44820 31168 44829
rect 32496 44863 32548 44872
rect 32496 44829 32505 44863
rect 32505 44829 32539 44863
rect 32539 44829 32548 44863
rect 32496 44820 32548 44829
rect 35440 44820 35492 44872
rect 20720 44752 20772 44804
rect 30012 44752 30064 44804
rect 30288 44795 30340 44804
rect 30288 44761 30297 44795
rect 30297 44761 30331 44795
rect 30331 44761 30340 44795
rect 30288 44752 30340 44761
rect 41420 44820 41472 44872
rect 41696 44863 41748 44872
rect 41696 44829 41705 44863
rect 41705 44829 41739 44863
rect 41739 44829 41748 44863
rect 41696 44820 41748 44829
rect 41788 44820 41840 44872
rect 44180 44888 44232 44940
rect 45744 44888 45796 44940
rect 47584 44931 47636 44940
rect 47584 44897 47593 44931
rect 47593 44897 47627 44931
rect 47627 44897 47636 44931
rect 47584 44888 47636 44897
rect 66260 44931 66312 44940
rect 66260 44897 66269 44931
rect 66269 44897 66303 44931
rect 66303 44897 66312 44931
rect 66260 44888 66312 44897
rect 68100 44931 68152 44940
rect 68100 44897 68109 44931
rect 68109 44897 68143 44931
rect 68143 44897 68152 44931
rect 68100 44888 68152 44897
rect 44364 44820 44416 44872
rect 45652 44820 45704 44872
rect 46204 44820 46256 44872
rect 21916 44684 21968 44736
rect 30932 44684 30984 44736
rect 34336 44684 34388 44736
rect 36176 44684 36228 44736
rect 43536 44752 43588 44804
rect 48320 44820 48372 44872
rect 51356 44820 51408 44872
rect 48412 44752 48464 44804
rect 66444 44795 66496 44804
rect 66444 44761 66453 44795
rect 66453 44761 66487 44795
rect 66487 44761 66496 44795
rect 66444 44752 66496 44761
rect 43812 44727 43864 44736
rect 43812 44693 43821 44727
rect 43821 44693 43855 44727
rect 43855 44693 43864 44727
rect 43812 44684 43864 44693
rect 44180 44684 44232 44736
rect 46664 44684 46716 44736
rect 47676 44684 47728 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 14556 44480 14608 44532
rect 12624 44387 12676 44396
rect 12624 44353 12633 44387
rect 12633 44353 12667 44387
rect 12667 44353 12676 44387
rect 12624 44344 12676 44353
rect 14740 44344 14792 44396
rect 15384 44387 15436 44396
rect 15384 44353 15393 44387
rect 15393 44353 15427 44387
rect 15427 44353 15436 44387
rect 15384 44344 15436 44353
rect 17040 44344 17092 44396
rect 20536 44480 20588 44532
rect 23296 44480 23348 44532
rect 29920 44480 29972 44532
rect 21916 44412 21968 44464
rect 21824 44344 21876 44396
rect 24032 44412 24084 44464
rect 30748 44455 30800 44464
rect 30748 44421 30757 44455
rect 30757 44421 30791 44455
rect 30791 44421 30800 44455
rect 30748 44412 30800 44421
rect 23572 44344 23624 44396
rect 25228 44387 25280 44396
rect 25228 44353 25237 44387
rect 25237 44353 25271 44387
rect 25271 44353 25280 44387
rect 25228 44344 25280 44353
rect 28908 44344 28960 44396
rect 34612 44480 34664 44532
rect 34704 44480 34756 44532
rect 17960 44319 18012 44328
rect 17960 44285 17969 44319
rect 17969 44285 18003 44319
rect 18003 44285 18012 44319
rect 17960 44276 18012 44285
rect 16764 44208 16816 44260
rect 18972 44319 19024 44328
rect 18972 44285 19006 44319
rect 19006 44285 19024 44319
rect 18972 44276 19024 44285
rect 19156 44319 19208 44328
rect 19156 44285 19165 44319
rect 19165 44285 19199 44319
rect 19199 44285 19208 44319
rect 19156 44276 19208 44285
rect 24032 44276 24084 44328
rect 34152 44344 34204 44396
rect 41696 44480 41748 44532
rect 44916 44480 44968 44532
rect 45836 44523 45888 44532
rect 45836 44489 45845 44523
rect 45845 44489 45879 44523
rect 45879 44489 45888 44523
rect 45836 44480 45888 44489
rect 47952 44523 48004 44532
rect 47952 44489 47961 44523
rect 47961 44489 47995 44523
rect 47995 44489 48004 44523
rect 47952 44480 48004 44489
rect 51356 44480 51408 44532
rect 66444 44480 66496 44532
rect 34796 44344 34848 44396
rect 36268 44412 36320 44464
rect 41052 44412 41104 44464
rect 41420 44344 41472 44396
rect 34520 44276 34572 44328
rect 34612 44276 34664 44328
rect 18328 44208 18380 44260
rect 42524 44344 42576 44396
rect 43812 44344 43864 44396
rect 45744 44344 45796 44396
rect 47676 44387 47728 44396
rect 43168 44319 43220 44328
rect 43168 44285 43177 44319
rect 43177 44285 43211 44319
rect 43211 44285 43220 44319
rect 43168 44276 43220 44285
rect 46204 44276 46256 44328
rect 47676 44353 47685 44387
rect 47685 44353 47719 44387
rect 47719 44353 47728 44387
rect 47676 44344 47728 44353
rect 47768 44387 47820 44396
rect 47768 44353 47777 44387
rect 47777 44353 47811 44387
rect 47811 44353 47820 44387
rect 48504 44387 48556 44396
rect 47768 44344 47820 44353
rect 48504 44353 48513 44387
rect 48513 44353 48547 44387
rect 48547 44353 48556 44387
rect 48504 44344 48556 44353
rect 48688 44344 48740 44396
rect 66628 44344 66680 44396
rect 42432 44208 42484 44260
rect 45652 44208 45704 44260
rect 12624 44183 12676 44192
rect 12624 44149 12633 44183
rect 12633 44149 12667 44183
rect 12667 44149 12676 44183
rect 12624 44140 12676 44149
rect 15200 44183 15252 44192
rect 15200 44149 15209 44183
rect 15209 44149 15243 44183
rect 15243 44149 15252 44183
rect 15200 44140 15252 44149
rect 16856 44140 16908 44192
rect 20996 44140 21048 44192
rect 22008 44140 22060 44192
rect 25044 44183 25096 44192
rect 25044 44149 25053 44183
rect 25053 44149 25087 44183
rect 25087 44149 25096 44183
rect 25044 44140 25096 44149
rect 27252 44140 27304 44192
rect 28356 44140 28408 44192
rect 30564 44140 30616 44192
rect 31208 44140 31260 44192
rect 32128 44183 32180 44192
rect 32128 44149 32137 44183
rect 32137 44149 32171 44183
rect 32171 44149 32180 44183
rect 32128 44140 32180 44149
rect 33784 44183 33836 44192
rect 33784 44149 33793 44183
rect 33793 44149 33827 44183
rect 33827 44149 33836 44183
rect 33784 44140 33836 44149
rect 36268 44140 36320 44192
rect 45560 44140 45612 44192
rect 48596 44183 48648 44192
rect 48596 44149 48605 44183
rect 48605 44149 48639 44183
rect 48639 44149 48648 44183
rect 48596 44140 48648 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 65654 44038 65706 44090
rect 65718 44038 65770 44090
rect 65782 44038 65834 44090
rect 65846 44038 65898 44090
rect 65910 44038 65962 44090
rect 20536 43936 20588 43988
rect 16580 43868 16632 43920
rect 16764 43868 16816 43920
rect 18328 43868 18380 43920
rect 19064 43868 19116 43920
rect 1860 43707 1912 43716
rect 1860 43673 1869 43707
rect 1869 43673 1903 43707
rect 1903 43673 1912 43707
rect 1860 43664 1912 43673
rect 13360 43775 13412 43784
rect 13360 43741 13369 43775
rect 13369 43741 13403 43775
rect 13403 43741 13412 43775
rect 14648 43775 14700 43784
rect 13360 43732 13412 43741
rect 14096 43664 14148 43716
rect 14648 43741 14657 43775
rect 14657 43741 14691 43775
rect 14691 43741 14700 43775
rect 14648 43732 14700 43741
rect 15200 43732 15252 43784
rect 15752 43664 15804 43716
rect 16856 43732 16908 43784
rect 25412 43868 25464 43920
rect 20996 43800 21048 43852
rect 21180 43732 21232 43784
rect 21364 43775 21416 43784
rect 21364 43741 21373 43775
rect 21373 43741 21407 43775
rect 21407 43741 21416 43775
rect 21364 43732 21416 43741
rect 20720 43664 20772 43716
rect 21824 43732 21876 43784
rect 29000 43936 29052 43988
rect 31208 43936 31260 43988
rect 34428 43936 34480 43988
rect 36360 43936 36412 43988
rect 28908 43868 28960 43920
rect 35808 43868 35860 43920
rect 40408 43936 40460 43988
rect 43168 43936 43220 43988
rect 44364 43979 44416 43988
rect 44364 43945 44373 43979
rect 44373 43945 44407 43979
rect 44407 43945 44416 43979
rect 44364 43936 44416 43945
rect 30932 43843 30984 43852
rect 22744 43775 22796 43784
rect 22744 43741 22753 43775
rect 22753 43741 22787 43775
rect 22787 43741 22796 43775
rect 22744 43732 22796 43741
rect 21916 43664 21968 43716
rect 24124 43732 24176 43784
rect 25044 43732 25096 43784
rect 13360 43596 13412 43648
rect 16764 43596 16816 43648
rect 20260 43596 20312 43648
rect 21088 43596 21140 43648
rect 21548 43596 21600 43648
rect 23020 43596 23072 43648
rect 24308 43596 24360 43648
rect 27160 43775 27212 43784
rect 27160 43741 27169 43775
rect 27169 43741 27203 43775
rect 27203 43741 27212 43775
rect 27160 43732 27212 43741
rect 26976 43596 27028 43648
rect 30932 43809 30941 43843
rect 30941 43809 30975 43843
rect 30975 43809 30984 43843
rect 30932 43800 30984 43809
rect 34520 43800 34572 43852
rect 36176 43800 36228 43852
rect 38660 43800 38712 43852
rect 38844 43800 38896 43852
rect 44916 43800 44968 43852
rect 45652 43843 45704 43852
rect 45652 43809 45661 43843
rect 45661 43809 45695 43843
rect 45695 43809 45704 43843
rect 45652 43800 45704 43809
rect 67916 43800 67968 43852
rect 28080 43775 28132 43784
rect 28080 43741 28089 43775
rect 28089 43741 28123 43775
rect 28123 43741 28132 43775
rect 28356 43775 28408 43784
rect 28080 43732 28132 43741
rect 28356 43741 28365 43775
rect 28365 43741 28399 43775
rect 28399 43741 28408 43775
rect 28356 43732 28408 43741
rect 29552 43707 29604 43716
rect 29552 43673 29561 43707
rect 29561 43673 29595 43707
rect 29595 43673 29604 43707
rect 29552 43664 29604 43673
rect 29920 43664 29972 43716
rect 32128 43732 32180 43784
rect 32772 43775 32824 43784
rect 32772 43741 32781 43775
rect 32781 43741 32815 43775
rect 32815 43741 32824 43775
rect 32772 43732 32824 43741
rect 33784 43732 33836 43784
rect 36268 43775 36320 43784
rect 36268 43741 36277 43775
rect 36277 43741 36311 43775
rect 36311 43741 36320 43775
rect 36268 43732 36320 43741
rect 37924 43775 37976 43784
rect 37924 43741 37933 43775
rect 37933 43741 37967 43775
rect 37967 43741 37976 43775
rect 37924 43732 37976 43741
rect 38108 43775 38160 43784
rect 38108 43741 38117 43775
rect 38117 43741 38151 43775
rect 38151 43741 38160 43775
rect 38108 43732 38160 43741
rect 38936 43732 38988 43784
rect 40500 43732 40552 43784
rect 42432 43775 42484 43784
rect 42432 43741 42441 43775
rect 42441 43741 42475 43775
rect 42475 43741 42484 43775
rect 42432 43732 42484 43741
rect 44180 43775 44232 43784
rect 44180 43741 44189 43775
rect 44189 43741 44223 43775
rect 44223 43741 44232 43775
rect 44180 43732 44232 43741
rect 46204 43732 46256 43784
rect 35992 43664 36044 43716
rect 38660 43707 38712 43716
rect 38660 43673 38669 43707
rect 38669 43673 38703 43707
rect 38703 43673 38712 43707
rect 38660 43664 38712 43673
rect 38844 43707 38896 43716
rect 38844 43673 38853 43707
rect 38853 43673 38887 43707
rect 38887 43673 38896 43707
rect 38844 43664 38896 43673
rect 42524 43664 42576 43716
rect 46388 43664 46440 43716
rect 48596 43732 48648 43784
rect 48320 43707 48372 43716
rect 48320 43673 48354 43707
rect 48354 43673 48372 43707
rect 66444 43707 66496 43716
rect 48320 43664 48372 43673
rect 66444 43673 66453 43707
rect 66453 43673 66487 43707
rect 66487 43673 66496 43707
rect 66444 43664 66496 43673
rect 68100 43707 68152 43716
rect 68100 43673 68109 43707
rect 68109 43673 68143 43707
rect 68143 43673 68152 43707
rect 68100 43664 68152 43673
rect 28816 43596 28868 43648
rect 30748 43596 30800 43648
rect 33600 43596 33652 43648
rect 38476 43596 38528 43648
rect 45652 43596 45704 43648
rect 47676 43596 47728 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 14648 43392 14700 43444
rect 15384 43392 15436 43444
rect 15752 43392 15804 43444
rect 17040 43435 17092 43444
rect 12624 43256 12676 43308
rect 12992 43299 13044 43308
rect 12992 43265 13026 43299
rect 13026 43265 13044 43299
rect 14556 43299 14608 43308
rect 12992 43256 13044 43265
rect 14556 43265 14565 43299
rect 14565 43265 14599 43299
rect 14599 43265 14608 43299
rect 14556 43256 14608 43265
rect 16580 43324 16632 43376
rect 15568 43256 15620 43308
rect 16764 43299 16816 43308
rect 16764 43265 16773 43299
rect 16773 43265 16807 43299
rect 16807 43265 16816 43299
rect 16764 43256 16816 43265
rect 17040 43401 17049 43435
rect 17049 43401 17083 43435
rect 17083 43401 17092 43435
rect 17040 43392 17092 43401
rect 19156 43392 19208 43444
rect 20444 43392 20496 43444
rect 20536 43392 20588 43444
rect 24124 43435 24176 43444
rect 24124 43401 24133 43435
rect 24133 43401 24167 43435
rect 24167 43401 24176 43435
rect 24124 43392 24176 43401
rect 25228 43392 25280 43444
rect 27160 43392 27212 43444
rect 29552 43392 29604 43444
rect 29644 43392 29696 43444
rect 30472 43392 30524 43444
rect 32772 43392 32824 43444
rect 34152 43435 34204 43444
rect 34152 43401 34161 43435
rect 34161 43401 34195 43435
rect 34195 43401 34204 43435
rect 34152 43392 34204 43401
rect 38844 43392 38896 43444
rect 39856 43392 39908 43444
rect 46388 43435 46440 43444
rect 46388 43401 46397 43435
rect 46397 43401 46431 43435
rect 46431 43401 46440 43435
rect 46388 43392 46440 43401
rect 48504 43392 48556 43444
rect 66444 43392 66496 43444
rect 25780 43324 25832 43376
rect 27252 43367 27304 43376
rect 27252 43333 27286 43367
rect 27286 43333 27304 43367
rect 27252 43324 27304 43333
rect 33600 43324 33652 43376
rect 33968 43367 34020 43376
rect 33968 43333 33993 43367
rect 33993 43333 34020 43367
rect 33968 43324 34020 43333
rect 34520 43324 34572 43376
rect 20260 43299 20312 43308
rect 20260 43265 20294 43299
rect 20294 43265 20312 43299
rect 22560 43299 22612 43308
rect 20260 43256 20312 43265
rect 22560 43265 22569 43299
rect 22569 43265 22603 43299
rect 22603 43265 22612 43299
rect 22560 43256 22612 43265
rect 24032 43299 24084 43308
rect 24032 43265 24041 43299
rect 24041 43265 24075 43299
rect 24075 43265 24084 43299
rect 24032 43256 24084 43265
rect 25412 43299 25464 43308
rect 25412 43265 25421 43299
rect 25421 43265 25455 43299
rect 25455 43265 25464 43299
rect 25412 43256 25464 43265
rect 26976 43299 27028 43308
rect 19340 43188 19392 43240
rect 20168 43231 20220 43240
rect 14096 43163 14148 43172
rect 14096 43129 14105 43163
rect 14105 43129 14139 43163
rect 14139 43129 14148 43163
rect 14096 43120 14148 43129
rect 18972 43120 19024 43172
rect 19064 43120 19116 43172
rect 20168 43197 20177 43231
rect 20177 43197 20211 43231
rect 20211 43197 20220 43231
rect 20168 43188 20220 43197
rect 20444 43231 20496 43240
rect 20444 43197 20453 43231
rect 20453 43197 20487 43231
rect 20487 43197 20496 43231
rect 20444 43188 20496 43197
rect 21180 43188 21232 43240
rect 25228 43188 25280 43240
rect 26976 43265 26985 43299
rect 26985 43265 27019 43299
rect 27019 43265 27028 43299
rect 26976 43256 27028 43265
rect 29000 43256 29052 43308
rect 21272 43120 21324 43172
rect 21640 43052 21692 43104
rect 29552 43256 29604 43308
rect 33876 43256 33928 43308
rect 37832 43256 37884 43308
rect 29460 43188 29512 43240
rect 30196 43231 30248 43240
rect 30196 43197 30230 43231
rect 30230 43197 30248 43231
rect 30196 43188 30248 43197
rect 30564 43188 30616 43240
rect 31024 43188 31076 43240
rect 38660 43324 38712 43376
rect 40500 43324 40552 43376
rect 39396 43256 39448 43308
rect 42524 43256 42576 43308
rect 45652 43299 45704 43308
rect 45652 43265 45661 43299
rect 45661 43265 45695 43299
rect 45695 43265 45704 43299
rect 45652 43256 45704 43265
rect 47676 43299 47728 43308
rect 38844 43231 38896 43240
rect 38844 43197 38853 43231
rect 38853 43197 38887 43231
rect 38887 43197 38896 43231
rect 38844 43188 38896 43197
rect 44180 43188 44232 43240
rect 47676 43265 47685 43299
rect 47685 43265 47719 43299
rect 47719 43265 47728 43299
rect 47676 43256 47728 43265
rect 47768 43299 47820 43308
rect 47768 43265 47777 43299
rect 47777 43265 47811 43299
rect 47811 43265 47820 43299
rect 47768 43256 47820 43265
rect 48688 43256 48740 43308
rect 66996 43256 67048 43308
rect 31760 43120 31812 43172
rect 35900 43120 35952 43172
rect 40960 43163 41012 43172
rect 40960 43129 40969 43163
rect 40969 43129 41003 43163
rect 41003 43129 41012 43163
rect 40960 43120 41012 43129
rect 30748 43052 30800 43104
rect 32956 43052 33008 43104
rect 34428 43052 34480 43104
rect 34520 43052 34572 43104
rect 41788 43095 41840 43104
rect 41788 43061 41797 43095
rect 41797 43061 41831 43095
rect 41831 43061 41840 43095
rect 41788 43052 41840 43061
rect 43812 43095 43864 43104
rect 43812 43061 43821 43095
rect 43821 43061 43855 43095
rect 43855 43061 43864 43095
rect 43812 43052 43864 43061
rect 48136 43052 48188 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 65654 42950 65706 43002
rect 65718 42950 65770 43002
rect 65782 42950 65834 43002
rect 65846 42950 65898 43002
rect 65910 42950 65962 43002
rect 12992 42848 13044 42900
rect 22744 42848 22796 42900
rect 31024 42848 31076 42900
rect 34428 42848 34480 42900
rect 38844 42848 38896 42900
rect 39948 42848 40000 42900
rect 32772 42823 32824 42832
rect 32772 42789 32781 42823
rect 32781 42789 32815 42823
rect 32815 42789 32824 42823
rect 32772 42780 32824 42789
rect 17960 42712 18012 42764
rect 21180 42712 21232 42764
rect 13360 42687 13412 42696
rect 13360 42653 13369 42687
rect 13369 42653 13403 42687
rect 13403 42653 13412 42687
rect 13360 42644 13412 42653
rect 14556 42644 14608 42696
rect 15752 42644 15804 42696
rect 16948 42687 17000 42696
rect 16948 42653 16957 42687
rect 16957 42653 16991 42687
rect 16991 42653 17000 42687
rect 16948 42644 17000 42653
rect 17500 42644 17552 42696
rect 25688 42712 25740 42764
rect 26056 42712 26108 42764
rect 28356 42712 28408 42764
rect 31760 42712 31812 42764
rect 36268 42712 36320 42764
rect 39856 42755 39908 42764
rect 21640 42687 21692 42696
rect 21640 42653 21649 42687
rect 21649 42653 21683 42687
rect 21683 42653 21692 42687
rect 21640 42644 21692 42653
rect 1860 42619 1912 42628
rect 1860 42585 1869 42619
rect 1869 42585 1903 42619
rect 1903 42585 1912 42619
rect 1860 42576 1912 42585
rect 18788 42576 18840 42628
rect 20996 42576 21048 42628
rect 22284 42576 22336 42628
rect 25044 42644 25096 42696
rect 26976 42644 27028 42696
rect 29552 42687 29604 42696
rect 29552 42653 29561 42687
rect 29561 42653 29595 42687
rect 29595 42653 29604 42687
rect 29552 42644 29604 42653
rect 24032 42576 24084 42628
rect 24492 42576 24544 42628
rect 1952 42551 2004 42560
rect 1952 42517 1961 42551
rect 1961 42517 1995 42551
rect 1995 42517 2004 42551
rect 1952 42508 2004 42517
rect 14740 42508 14792 42560
rect 15476 42551 15528 42560
rect 15476 42517 15485 42551
rect 15485 42517 15519 42551
rect 15519 42517 15528 42551
rect 15476 42508 15528 42517
rect 16948 42508 17000 42560
rect 17960 42551 18012 42560
rect 17960 42517 17969 42551
rect 17969 42517 18003 42551
rect 18003 42517 18012 42551
rect 17960 42508 18012 42517
rect 21548 42551 21600 42560
rect 21548 42517 21557 42551
rect 21557 42517 21591 42551
rect 21591 42517 21600 42551
rect 21548 42508 21600 42517
rect 23664 42508 23716 42560
rect 29736 42576 29788 42628
rect 30748 42644 30800 42696
rect 32772 42644 32824 42696
rect 34152 42644 34204 42696
rect 37372 42644 37424 42696
rect 37924 42644 37976 42696
rect 39856 42721 39865 42755
rect 39865 42721 39899 42755
rect 39899 42721 39908 42755
rect 39856 42712 39908 42721
rect 46572 42712 46624 42764
rect 67916 42755 67968 42764
rect 67916 42721 67925 42755
rect 67925 42721 67959 42755
rect 67959 42721 67968 42755
rect 67916 42712 67968 42721
rect 29920 42576 29972 42628
rect 24952 42508 25004 42560
rect 30196 42508 30248 42560
rect 31116 42508 31168 42560
rect 31760 42551 31812 42560
rect 31760 42517 31769 42551
rect 31769 42517 31803 42551
rect 31803 42517 31812 42551
rect 32496 42576 32548 42628
rect 33784 42619 33836 42628
rect 33784 42585 33793 42619
rect 33793 42585 33827 42619
rect 33827 42585 33836 42619
rect 33784 42576 33836 42585
rect 35440 42576 35492 42628
rect 37648 42576 37700 42628
rect 38016 42576 38068 42628
rect 40132 42644 40184 42696
rect 40316 42644 40368 42696
rect 41788 42644 41840 42696
rect 41880 42644 41932 42696
rect 43352 42644 43404 42696
rect 48136 42687 48188 42696
rect 48136 42653 48145 42687
rect 48145 42653 48179 42687
rect 48179 42653 48188 42687
rect 48136 42644 48188 42653
rect 65800 42644 65852 42696
rect 44088 42619 44140 42628
rect 31760 42508 31812 42517
rect 33968 42551 34020 42560
rect 33968 42517 33993 42551
rect 33993 42517 34020 42551
rect 33968 42508 34020 42517
rect 35716 42508 35768 42560
rect 36084 42551 36136 42560
rect 36084 42517 36093 42551
rect 36093 42517 36127 42551
rect 36127 42517 36136 42551
rect 36084 42508 36136 42517
rect 37832 42508 37884 42560
rect 39764 42508 39816 42560
rect 41328 42508 41380 42560
rect 44088 42585 44097 42619
rect 44097 42585 44131 42619
rect 44131 42585 44140 42619
rect 44088 42576 44140 42585
rect 45284 42576 45336 42628
rect 45008 42551 45060 42560
rect 45008 42517 45017 42551
rect 45017 42517 45051 42551
rect 45051 42517 45060 42551
rect 45008 42508 45060 42517
rect 48320 42508 48372 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 1952 42304 2004 42356
rect 15476 42236 15528 42288
rect 14740 42211 14792 42220
rect 14740 42177 14749 42211
rect 14749 42177 14783 42211
rect 14783 42177 14792 42211
rect 14740 42168 14792 42177
rect 16948 42211 17000 42220
rect 16948 42177 16957 42211
rect 16957 42177 16991 42211
rect 16991 42177 17000 42211
rect 16948 42168 17000 42177
rect 17224 42211 17276 42220
rect 17224 42177 17258 42211
rect 17258 42177 17276 42211
rect 18052 42304 18104 42356
rect 18420 42304 18472 42356
rect 25044 42304 25096 42356
rect 25872 42304 25924 42356
rect 28356 42347 28408 42356
rect 28356 42313 28365 42347
rect 28365 42313 28399 42347
rect 28399 42313 28408 42347
rect 28356 42304 28408 42313
rect 29736 42304 29788 42356
rect 31024 42304 31076 42356
rect 32128 42304 32180 42356
rect 34152 42347 34204 42356
rect 17500 42236 17552 42288
rect 18788 42211 18840 42220
rect 17224 42168 17276 42177
rect 18788 42177 18797 42211
rect 18797 42177 18831 42211
rect 18831 42177 18840 42211
rect 18788 42168 18840 42177
rect 19340 42168 19392 42220
rect 19616 42211 19668 42220
rect 19616 42177 19625 42211
rect 19625 42177 19659 42211
rect 19659 42177 19668 42211
rect 19616 42168 19668 42177
rect 30748 42236 30800 42288
rect 31760 42236 31812 42288
rect 34152 42313 34161 42347
rect 34161 42313 34195 42347
rect 34195 42313 34204 42347
rect 34152 42304 34204 42313
rect 35440 42347 35492 42356
rect 35440 42313 35449 42347
rect 35449 42313 35483 42347
rect 35483 42313 35492 42347
rect 35440 42304 35492 42313
rect 35532 42304 35584 42356
rect 67088 42304 67140 42356
rect 20996 42168 21048 42220
rect 23388 42211 23440 42220
rect 22100 42100 22152 42152
rect 16120 42007 16172 42016
rect 16120 41973 16129 42007
rect 16129 41973 16163 42007
rect 16163 41973 16172 42007
rect 20168 42032 20220 42084
rect 23388 42177 23397 42211
rect 23397 42177 23431 42211
rect 23431 42177 23440 42211
rect 23388 42168 23440 42177
rect 24952 42211 25004 42220
rect 23572 42100 23624 42152
rect 24216 42100 24268 42152
rect 24308 42032 24360 42084
rect 24952 42177 24961 42211
rect 24961 42177 24995 42211
rect 24995 42177 25004 42211
rect 24952 42168 25004 42177
rect 25228 42168 25280 42220
rect 25412 42168 25464 42220
rect 26148 42211 26200 42220
rect 26148 42177 26157 42211
rect 26157 42177 26191 42211
rect 26191 42177 26200 42211
rect 26148 42168 26200 42177
rect 26976 42211 27028 42220
rect 26976 42177 26985 42211
rect 26985 42177 27019 42211
rect 27019 42177 27028 42211
rect 26976 42168 27028 42177
rect 25964 42143 26016 42152
rect 25964 42109 25973 42143
rect 25973 42109 26007 42143
rect 26007 42109 26016 42143
rect 25964 42100 26016 42109
rect 27528 42168 27580 42220
rect 28632 42168 28684 42220
rect 29092 42211 29144 42220
rect 29092 42177 29101 42211
rect 29101 42177 29135 42211
rect 29135 42177 29144 42211
rect 29092 42168 29144 42177
rect 31116 42168 31168 42220
rect 32772 42168 32824 42220
rect 32956 42168 33008 42220
rect 33968 42211 34020 42220
rect 29184 42100 29236 42152
rect 29368 42100 29420 42152
rect 16120 41964 16172 41973
rect 19248 41964 19300 42016
rect 19984 41964 20036 42016
rect 24032 42007 24084 42016
rect 24032 41973 24041 42007
rect 24041 41973 24075 42007
rect 24075 41973 24084 42007
rect 24032 41964 24084 41973
rect 24584 41964 24636 42016
rect 25872 42007 25924 42016
rect 25872 41973 25881 42007
rect 25881 41973 25915 42007
rect 25915 41973 25924 42007
rect 25872 41964 25924 41973
rect 26056 41964 26108 42016
rect 30104 42032 30156 42084
rect 33968 42177 33977 42211
rect 33977 42177 34011 42211
rect 34011 42177 34020 42211
rect 33968 42168 34020 42177
rect 37924 42236 37976 42288
rect 41880 42236 41932 42288
rect 43352 42279 43404 42288
rect 43352 42245 43361 42279
rect 43361 42245 43395 42279
rect 43395 42245 43404 42279
rect 43352 42236 43404 42245
rect 45008 42236 45060 42288
rect 35532 42168 35584 42220
rect 35716 42168 35768 42220
rect 35992 42168 36044 42220
rect 36544 42211 36596 42220
rect 36544 42177 36553 42211
rect 36553 42177 36587 42211
rect 36587 42177 36596 42211
rect 36544 42168 36596 42177
rect 33416 42100 33468 42152
rect 33784 42100 33836 42152
rect 36084 42100 36136 42152
rect 37372 42168 37424 42220
rect 39580 42168 39632 42220
rect 39764 42211 39816 42220
rect 39764 42177 39773 42211
rect 39773 42177 39807 42211
rect 39807 42177 39816 42211
rect 39764 42168 39816 42177
rect 41328 42211 41380 42220
rect 41328 42177 41337 42211
rect 41337 42177 41371 42211
rect 41371 42177 41380 42211
rect 41328 42168 41380 42177
rect 41696 42168 41748 42220
rect 43628 42168 43680 42220
rect 43812 42211 43864 42220
rect 43812 42177 43821 42211
rect 43821 42177 43855 42211
rect 43855 42177 43864 42211
rect 43812 42168 43864 42177
rect 65800 42211 65852 42220
rect 65800 42177 65809 42211
rect 65809 42177 65843 42211
rect 65843 42177 65852 42211
rect 65800 42168 65852 42177
rect 39028 42100 39080 42152
rect 42432 42100 42484 42152
rect 48596 42143 48648 42152
rect 38936 42032 38988 42084
rect 39212 42032 39264 42084
rect 39396 42032 39448 42084
rect 43168 42032 43220 42084
rect 28908 42007 28960 42016
rect 28908 41973 28917 42007
rect 28917 41973 28951 42007
rect 28951 41973 28960 42007
rect 28908 41964 28960 41973
rect 29184 41964 29236 42016
rect 32128 41964 32180 42016
rect 32496 41964 32548 42016
rect 34796 41964 34848 42016
rect 37648 42007 37700 42016
rect 37648 41973 37657 42007
rect 37657 41973 37691 42007
rect 37691 41973 37700 42007
rect 37648 41964 37700 41973
rect 38844 41964 38896 42016
rect 48596 42109 48605 42143
rect 48605 42109 48639 42143
rect 48639 42109 48648 42143
rect 48596 42100 48648 42109
rect 49424 42100 49476 42152
rect 64880 42100 64932 42152
rect 65984 42143 66036 42152
rect 65984 42109 65993 42143
rect 65993 42109 66027 42143
rect 66027 42109 66036 42143
rect 65984 42100 66036 42109
rect 67548 42143 67600 42152
rect 67548 42109 67557 42143
rect 67557 42109 67591 42143
rect 67591 42109 67600 42143
rect 67548 42100 67600 42109
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 65654 41862 65706 41914
rect 65718 41862 65770 41914
rect 65782 41862 65834 41914
rect 65846 41862 65898 41914
rect 65910 41862 65962 41914
rect 15752 41803 15804 41812
rect 15752 41769 15761 41803
rect 15761 41769 15795 41803
rect 15795 41769 15804 41803
rect 15752 41760 15804 41769
rect 14832 41692 14884 41744
rect 16120 41624 16172 41676
rect 18420 41692 18472 41744
rect 15568 41599 15620 41608
rect 15568 41565 15577 41599
rect 15577 41565 15611 41599
rect 15611 41565 15620 41599
rect 15568 41556 15620 41565
rect 17592 41599 17644 41608
rect 17592 41565 17601 41599
rect 17601 41565 17635 41599
rect 17635 41565 17644 41599
rect 17592 41556 17644 41565
rect 19616 41760 19668 41812
rect 19248 41667 19300 41676
rect 19248 41633 19257 41667
rect 19257 41633 19291 41667
rect 19291 41633 19300 41667
rect 19248 41624 19300 41633
rect 23664 41760 23716 41812
rect 24492 41760 24544 41812
rect 25780 41803 25832 41812
rect 25780 41769 25789 41803
rect 25789 41769 25823 41803
rect 25823 41769 25832 41803
rect 25780 41760 25832 41769
rect 26332 41760 26384 41812
rect 26516 41760 26568 41812
rect 27528 41760 27580 41812
rect 58716 41760 58768 41812
rect 65984 41760 66036 41812
rect 29000 41735 29052 41744
rect 29000 41701 29009 41735
rect 29009 41701 29043 41735
rect 29043 41701 29052 41735
rect 29000 41692 29052 41701
rect 29460 41692 29512 41744
rect 31024 41692 31076 41744
rect 37280 41692 37332 41744
rect 39028 41692 39080 41744
rect 22100 41624 22152 41676
rect 21180 41556 21232 41608
rect 23572 41556 23624 41608
rect 24584 41599 24636 41608
rect 24584 41565 24593 41599
rect 24593 41565 24627 41599
rect 24627 41565 24636 41599
rect 24584 41556 24636 41565
rect 17684 41488 17736 41540
rect 19432 41420 19484 41472
rect 21824 41488 21876 41540
rect 21916 41420 21968 41472
rect 23112 41420 23164 41472
rect 23388 41420 23440 41472
rect 26332 41556 26384 41608
rect 27712 41556 27764 41608
rect 28172 41556 28224 41608
rect 28908 41488 28960 41540
rect 29920 41599 29972 41608
rect 29920 41565 29929 41599
rect 29929 41565 29963 41599
rect 29963 41565 29972 41599
rect 38384 41624 38436 41676
rect 29920 41556 29972 41565
rect 32772 41556 32824 41608
rect 33968 41556 34020 41608
rect 35440 41599 35492 41608
rect 35440 41565 35449 41599
rect 35449 41565 35483 41599
rect 35483 41565 35492 41599
rect 35440 41556 35492 41565
rect 35532 41556 35584 41608
rect 38292 41556 38344 41608
rect 38660 41556 38712 41608
rect 30656 41488 30708 41540
rect 34796 41488 34848 41540
rect 36544 41531 36596 41540
rect 36544 41497 36553 41531
rect 36553 41497 36587 41531
rect 36587 41497 36596 41531
rect 36544 41488 36596 41497
rect 37280 41488 37332 41540
rect 38108 41488 38160 41540
rect 38844 41599 38896 41608
rect 38844 41565 38858 41599
rect 38858 41565 38892 41599
rect 38892 41565 38896 41599
rect 38844 41556 38896 41565
rect 39580 41624 39632 41676
rect 42248 41667 42300 41676
rect 42248 41633 42280 41667
rect 42280 41633 42300 41667
rect 42248 41624 42300 41633
rect 42432 41667 42484 41676
rect 42432 41633 42441 41667
rect 42441 41633 42475 41667
rect 42475 41633 42484 41667
rect 42432 41624 42484 41633
rect 41328 41556 41380 41608
rect 42340 41599 42392 41608
rect 38936 41488 38988 41540
rect 29184 41420 29236 41472
rect 31300 41463 31352 41472
rect 31300 41429 31309 41463
rect 31309 41429 31343 41463
rect 31343 41429 31352 41463
rect 31300 41420 31352 41429
rect 32772 41420 32824 41472
rect 35256 41463 35308 41472
rect 35256 41429 35265 41463
rect 35265 41429 35299 41463
rect 35299 41429 35308 41463
rect 35256 41420 35308 41429
rect 37464 41420 37516 41472
rect 37740 41420 37792 41472
rect 39028 41420 39080 41472
rect 41512 41488 41564 41540
rect 42340 41565 42349 41599
rect 42349 41565 42383 41599
rect 42383 41565 42392 41599
rect 42340 41556 42392 41565
rect 45376 41624 45428 41676
rect 43168 41599 43220 41608
rect 43168 41565 43177 41599
rect 43177 41565 43211 41599
rect 43211 41565 43220 41599
rect 43168 41556 43220 41565
rect 45468 41599 45520 41608
rect 45468 41565 45477 41599
rect 45477 41565 45511 41599
rect 45511 41565 45520 41599
rect 45468 41556 45520 41565
rect 45744 41556 45796 41608
rect 46296 41692 46348 41744
rect 49424 41735 49476 41744
rect 49424 41701 49433 41735
rect 49433 41701 49467 41735
rect 49467 41701 49476 41735
rect 49424 41692 49476 41701
rect 48780 41556 48832 41608
rect 66996 41556 67048 41608
rect 42892 41488 42944 41540
rect 41972 41463 42024 41472
rect 41972 41429 41981 41463
rect 41981 41429 42015 41463
rect 42015 41429 42024 41463
rect 41972 41420 42024 41429
rect 42340 41420 42392 41472
rect 42800 41420 42852 41472
rect 46664 41488 46716 41540
rect 45652 41420 45704 41472
rect 48596 41420 48648 41472
rect 48872 41420 48924 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 17224 41216 17276 41268
rect 19432 41259 19484 41268
rect 19432 41225 19441 41259
rect 19441 41225 19475 41259
rect 19475 41225 19484 41259
rect 19432 41216 19484 41225
rect 21824 41259 21876 41268
rect 21824 41225 21833 41259
rect 21833 41225 21867 41259
rect 21867 41225 21876 41259
rect 21824 41216 21876 41225
rect 23296 41216 23348 41268
rect 23480 41148 23532 41200
rect 24032 41148 24084 41200
rect 27712 41191 27764 41200
rect 17960 41080 18012 41132
rect 19984 41080 20036 41132
rect 19248 41012 19300 41064
rect 21916 41012 21968 41064
rect 22192 41089 22201 41116
rect 22201 41089 22235 41116
rect 22235 41089 22244 41116
rect 22192 41064 22244 41089
rect 22284 41123 22336 41132
rect 22284 41089 22293 41123
rect 22293 41089 22327 41123
rect 22327 41089 22336 41123
rect 22284 41080 22336 41089
rect 23664 41080 23716 41132
rect 24952 41123 25004 41132
rect 24952 41089 24961 41123
rect 24961 41089 24995 41123
rect 24995 41089 25004 41123
rect 24952 41080 25004 41089
rect 27712 41157 27721 41191
rect 27721 41157 27755 41191
rect 27755 41157 27764 41191
rect 27712 41148 27764 41157
rect 29092 41216 29144 41268
rect 29920 41216 29972 41268
rect 30656 41259 30708 41268
rect 30656 41225 30665 41259
rect 30665 41225 30699 41259
rect 30699 41225 30708 41259
rect 30656 41216 30708 41225
rect 42340 41216 42392 41268
rect 45744 41216 45796 41268
rect 35256 41148 35308 41200
rect 37556 41148 37608 41200
rect 39028 41148 39080 41200
rect 42524 41148 42576 41200
rect 42892 41148 42944 41200
rect 45376 41148 45428 41200
rect 28448 41123 28500 41132
rect 24400 40944 24452 40996
rect 27252 40944 27304 40996
rect 28448 41089 28457 41123
rect 28457 41089 28491 41123
rect 28491 41089 28500 41123
rect 28448 41080 28500 41089
rect 28264 41012 28316 41064
rect 29092 41080 29144 41132
rect 32496 41123 32548 41132
rect 32496 41089 32505 41123
rect 32505 41089 32539 41123
rect 32539 41089 32548 41123
rect 32496 41080 32548 41089
rect 32680 41123 32732 41132
rect 32680 41089 32689 41123
rect 32689 41089 32723 41123
rect 32723 41089 32732 41123
rect 32680 41080 32732 41089
rect 34428 41080 34480 41132
rect 37280 41123 37332 41132
rect 37280 41089 37289 41123
rect 37289 41089 37323 41123
rect 37323 41089 37332 41123
rect 37280 41080 37332 41089
rect 37464 41123 37516 41132
rect 37464 41089 37473 41123
rect 37473 41089 37507 41123
rect 37507 41089 37516 41123
rect 37464 41080 37516 41089
rect 37740 41080 37792 41132
rect 37832 41080 37884 41132
rect 38108 41123 38160 41132
rect 38108 41089 38117 41123
rect 38117 41089 38151 41123
rect 38151 41089 38160 41123
rect 38108 41080 38160 41089
rect 38384 41080 38436 41132
rect 31300 41012 31352 41064
rect 33508 41055 33560 41064
rect 33508 41021 33542 41055
rect 33542 41021 33560 41055
rect 33508 41012 33560 41021
rect 34520 41012 34572 41064
rect 38660 41012 38712 41064
rect 29092 40944 29144 40996
rect 24676 40876 24728 40928
rect 25872 40876 25924 40928
rect 26056 40876 26108 40928
rect 28448 40876 28500 40928
rect 29000 40876 29052 40928
rect 37556 40944 37608 40996
rect 38936 40944 38988 40996
rect 33876 40876 33928 40928
rect 35532 40876 35584 40928
rect 35624 40876 35676 40928
rect 37648 40919 37700 40928
rect 37648 40885 37657 40919
rect 37657 40885 37691 40919
rect 37691 40885 37700 40919
rect 37648 40876 37700 40885
rect 38384 40876 38436 40928
rect 40132 41012 40184 41064
rect 41512 41012 41564 41064
rect 42616 41055 42668 41064
rect 42616 41021 42625 41055
rect 42625 41021 42659 41055
rect 42659 41021 42668 41055
rect 42616 41012 42668 41021
rect 42800 41055 42852 41064
rect 42800 41021 42809 41055
rect 42809 41021 42843 41055
rect 42843 41021 42852 41055
rect 42800 41012 42852 41021
rect 42892 41055 42944 41064
rect 42892 41021 42901 41055
rect 42901 41021 42935 41055
rect 42935 41021 42944 41055
rect 43904 41080 43956 41132
rect 45928 41080 45980 41132
rect 46296 41148 46348 41200
rect 48872 41191 48924 41200
rect 48872 41157 48881 41191
rect 48881 41157 48915 41191
rect 48915 41157 48924 41191
rect 48872 41148 48924 41157
rect 42892 41012 42944 41021
rect 40960 40944 41012 40996
rect 67272 41080 67324 41132
rect 46296 41012 46348 41064
rect 48044 41012 48096 41064
rect 40316 40919 40368 40928
rect 40316 40885 40325 40919
rect 40325 40885 40359 40919
rect 40359 40885 40368 40919
rect 40316 40876 40368 40885
rect 41972 40876 42024 40928
rect 46388 40944 46440 40996
rect 60740 41012 60792 41064
rect 43628 40919 43680 40928
rect 43628 40885 43637 40919
rect 43637 40885 43671 40919
rect 43671 40885 43680 40919
rect 43628 40876 43680 40885
rect 44180 40919 44232 40928
rect 44180 40885 44189 40919
rect 44189 40885 44223 40919
rect 44223 40885 44232 40919
rect 44180 40876 44232 40885
rect 45744 40919 45796 40928
rect 45744 40885 45753 40919
rect 45753 40885 45787 40919
rect 45787 40885 45796 40919
rect 45744 40876 45796 40885
rect 66260 40876 66312 40928
rect 67088 40876 67140 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 65654 40774 65706 40826
rect 65718 40774 65770 40826
rect 65782 40774 65834 40826
rect 65846 40774 65898 40826
rect 65910 40774 65962 40826
rect 3240 40400 3292 40452
rect 19248 40579 19300 40588
rect 19248 40545 19257 40579
rect 19257 40545 19291 40579
rect 19291 40545 19300 40579
rect 19248 40536 19300 40545
rect 21272 40468 21324 40520
rect 22192 40672 22244 40724
rect 22744 40672 22796 40724
rect 22008 40604 22060 40656
rect 34520 40672 34572 40724
rect 34796 40672 34848 40724
rect 35348 40715 35400 40724
rect 35348 40681 35357 40715
rect 35357 40681 35391 40715
rect 35391 40681 35400 40715
rect 35348 40672 35400 40681
rect 35440 40672 35492 40724
rect 37832 40672 37884 40724
rect 42616 40672 42668 40724
rect 43904 40715 43956 40724
rect 43904 40681 43913 40715
rect 43913 40681 43947 40715
rect 43947 40681 43956 40715
rect 43904 40672 43956 40681
rect 48044 40715 48096 40724
rect 48044 40681 48053 40715
rect 48053 40681 48087 40715
rect 48087 40681 48096 40715
rect 48044 40672 48096 40681
rect 23664 40536 23716 40588
rect 24400 40579 24452 40588
rect 24400 40545 24409 40579
rect 24409 40545 24443 40579
rect 24443 40545 24452 40579
rect 24400 40536 24452 40545
rect 37556 40604 37608 40656
rect 37648 40604 37700 40656
rect 28080 40579 28132 40588
rect 28080 40545 28089 40579
rect 28089 40545 28123 40579
rect 28123 40545 28132 40579
rect 28080 40536 28132 40545
rect 29276 40536 29328 40588
rect 37280 40536 37332 40588
rect 38476 40579 38528 40588
rect 38476 40545 38485 40579
rect 38485 40545 38519 40579
rect 38519 40545 38528 40579
rect 38476 40536 38528 40545
rect 41420 40604 41472 40656
rect 39028 40536 39080 40588
rect 42340 40536 42392 40588
rect 45008 40536 45060 40588
rect 46664 40579 46716 40588
rect 23296 40468 23348 40520
rect 24676 40511 24728 40520
rect 24676 40477 24710 40511
rect 24710 40477 24728 40511
rect 24676 40468 24728 40477
rect 26240 40511 26292 40520
rect 26240 40477 26249 40511
rect 26249 40477 26283 40511
rect 26283 40477 26292 40511
rect 26240 40468 26292 40477
rect 28264 40511 28316 40520
rect 28264 40477 28273 40511
rect 28273 40477 28307 40511
rect 28307 40477 28316 40511
rect 28264 40468 28316 40477
rect 29092 40468 29144 40520
rect 33048 40468 33100 40520
rect 26976 40400 27028 40452
rect 19984 40332 20036 40384
rect 21548 40375 21600 40384
rect 21548 40341 21557 40375
rect 21557 40341 21591 40375
rect 21591 40341 21600 40375
rect 21548 40332 21600 40341
rect 23388 40375 23440 40384
rect 23388 40341 23397 40375
rect 23397 40341 23431 40375
rect 23431 40341 23440 40375
rect 23388 40332 23440 40341
rect 25136 40332 25188 40384
rect 33508 40400 33560 40452
rect 35164 40443 35216 40452
rect 35164 40409 35173 40443
rect 35173 40409 35207 40443
rect 35207 40409 35216 40443
rect 35164 40400 35216 40409
rect 35624 40400 35676 40452
rect 37372 40468 37424 40520
rect 39120 40468 39172 40520
rect 39396 40468 39448 40520
rect 37740 40400 37792 40452
rect 38660 40400 38712 40452
rect 39764 40400 39816 40452
rect 42524 40443 42576 40452
rect 42524 40409 42533 40443
rect 42533 40409 42567 40443
rect 42567 40409 42576 40443
rect 42524 40400 42576 40409
rect 43720 40511 43772 40520
rect 43720 40477 43729 40511
rect 43729 40477 43763 40511
rect 43763 40477 43772 40511
rect 46664 40545 46673 40579
rect 46673 40545 46707 40579
rect 46707 40545 46716 40579
rect 46664 40536 46716 40545
rect 66260 40579 66312 40588
rect 66260 40545 66269 40579
rect 66269 40545 66303 40579
rect 66303 40545 66312 40579
rect 66260 40536 66312 40545
rect 67088 40536 67140 40588
rect 68100 40579 68152 40588
rect 68100 40545 68109 40579
rect 68109 40545 68143 40579
rect 68143 40545 68152 40579
rect 68100 40536 68152 40545
rect 43720 40468 43772 40477
rect 45744 40468 45796 40520
rect 48780 40511 48832 40520
rect 48780 40477 48789 40511
rect 48789 40477 48823 40511
rect 48823 40477 48832 40511
rect 48780 40468 48832 40477
rect 45192 40400 45244 40452
rect 28448 40375 28500 40384
rect 28448 40341 28457 40375
rect 28457 40341 28491 40375
rect 28491 40341 28500 40375
rect 28448 40332 28500 40341
rect 29276 40332 29328 40384
rect 34704 40332 34756 40384
rect 35348 40375 35400 40384
rect 35348 40341 35373 40375
rect 35373 40341 35400 40375
rect 35348 40332 35400 40341
rect 38016 40332 38068 40384
rect 38752 40332 38804 40384
rect 46112 40332 46164 40384
rect 48964 40332 49016 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 22468 40128 22520 40180
rect 24952 40128 25004 40180
rect 26240 40128 26292 40180
rect 26976 40171 27028 40180
rect 26976 40137 26985 40171
rect 26985 40137 27019 40171
rect 27019 40137 27028 40171
rect 26976 40128 27028 40137
rect 19984 39992 20036 40044
rect 21548 39992 21600 40044
rect 23388 40060 23440 40112
rect 22836 39992 22888 40044
rect 25136 40035 25188 40044
rect 25136 40001 25145 40035
rect 25145 40001 25179 40035
rect 25179 40001 25188 40035
rect 25136 39992 25188 40001
rect 25228 40035 25280 40044
rect 25228 40001 25237 40035
rect 25237 40001 25271 40035
rect 25271 40001 25280 40035
rect 26332 40035 26384 40044
rect 25228 39992 25280 40001
rect 26332 40001 26341 40035
rect 26341 40001 26375 40035
rect 26375 40001 26384 40035
rect 26332 39992 26384 40001
rect 28448 40060 28500 40112
rect 28264 40035 28316 40044
rect 28264 40001 28273 40035
rect 28273 40001 28307 40035
rect 28307 40001 28316 40035
rect 28264 39992 28316 40001
rect 29276 40035 29328 40044
rect 29276 40001 29285 40035
rect 29285 40001 29319 40035
rect 29319 40001 29328 40035
rect 29276 39992 29328 40001
rect 30472 39992 30524 40044
rect 32312 40035 32364 40044
rect 32312 40001 32321 40035
rect 32321 40001 32355 40035
rect 32355 40001 32364 40035
rect 32312 39992 32364 40001
rect 33232 40035 33284 40044
rect 33232 40001 33241 40035
rect 33241 40001 33275 40035
rect 33275 40001 33284 40035
rect 33232 39992 33284 40001
rect 35164 40128 35216 40180
rect 38108 40128 38160 40180
rect 44364 40128 44416 40180
rect 45192 40171 45244 40180
rect 45192 40137 45201 40171
rect 45201 40137 45235 40171
rect 45235 40137 45244 40171
rect 45192 40128 45244 40137
rect 46296 40128 46348 40180
rect 38200 40103 38252 40112
rect 38200 40069 38209 40103
rect 38209 40069 38243 40103
rect 38243 40069 38252 40103
rect 38200 40060 38252 40069
rect 39212 40060 39264 40112
rect 39580 40060 39632 40112
rect 41420 40060 41472 40112
rect 42524 40103 42576 40112
rect 42524 40069 42533 40103
rect 42533 40069 42567 40103
rect 42567 40069 42576 40103
rect 42524 40060 42576 40069
rect 43352 40060 43404 40112
rect 44180 40060 44232 40112
rect 48136 40060 48188 40112
rect 48964 40103 49016 40112
rect 48964 40069 48973 40103
rect 48973 40069 49007 40103
rect 49007 40069 49016 40103
rect 48964 40060 49016 40069
rect 66076 40060 66128 40112
rect 67272 40103 67324 40112
rect 67272 40069 67281 40103
rect 67281 40069 67315 40103
rect 67315 40069 67324 40103
rect 67272 40060 67324 40069
rect 37832 39992 37884 40044
rect 40500 39992 40552 40044
rect 43628 39992 43680 40044
rect 46296 39992 46348 40044
rect 27804 39924 27856 39976
rect 32680 39924 32732 39976
rect 34244 39967 34296 39976
rect 34244 39933 34278 39967
rect 34278 39933 34296 39967
rect 34244 39924 34296 39933
rect 34796 39924 34848 39976
rect 39948 39967 40000 39976
rect 39948 39933 39957 39967
rect 39957 39933 39991 39967
rect 39991 39933 40000 39967
rect 39948 39924 40000 39933
rect 1400 39788 1452 39840
rect 21272 39831 21324 39840
rect 21272 39797 21281 39831
rect 21281 39797 21315 39831
rect 21315 39797 21324 39831
rect 21272 39788 21324 39797
rect 30564 39788 30616 39840
rect 33232 39856 33284 39908
rect 33600 39856 33652 39908
rect 33876 39899 33928 39908
rect 33876 39865 33885 39899
rect 33885 39865 33919 39899
rect 33919 39865 33928 39899
rect 33876 39856 33928 39865
rect 37924 39856 37976 39908
rect 38384 39899 38436 39908
rect 38384 39865 38393 39899
rect 38393 39865 38427 39899
rect 38427 39865 38436 39899
rect 38384 39856 38436 39865
rect 45376 39856 45428 39908
rect 46572 40038 46624 40044
rect 46572 40004 46581 40038
rect 46581 40004 46615 40038
rect 46615 40004 46624 40038
rect 46572 39992 46624 40004
rect 46756 40035 46808 40044
rect 46756 40001 46765 40035
rect 46765 40001 46799 40035
rect 46799 40001 46808 40035
rect 46756 39992 46808 40001
rect 31392 39831 31444 39840
rect 31392 39797 31401 39831
rect 31401 39797 31435 39831
rect 31435 39797 31444 39831
rect 31392 39788 31444 39797
rect 37648 39831 37700 39840
rect 37648 39797 37657 39831
rect 37657 39797 37691 39831
rect 37691 39797 37700 39831
rect 37648 39788 37700 39797
rect 39120 39831 39172 39840
rect 39120 39797 39129 39831
rect 39129 39797 39163 39831
rect 39163 39797 39172 39831
rect 39120 39788 39172 39797
rect 41052 39788 41104 39840
rect 42616 39788 42668 39840
rect 46848 39788 46900 39840
rect 67364 39831 67416 39840
rect 67364 39797 67373 39831
rect 67373 39797 67407 39831
rect 67407 39797 67416 39831
rect 67364 39788 67416 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 65654 39686 65706 39738
rect 65718 39686 65770 39738
rect 65782 39686 65834 39738
rect 65846 39686 65898 39738
rect 65910 39686 65962 39738
rect 25780 39627 25832 39636
rect 25780 39593 25789 39627
rect 25789 39593 25823 39627
rect 25823 39593 25832 39627
rect 25780 39584 25832 39593
rect 26148 39584 26200 39636
rect 26332 39584 26384 39636
rect 27252 39584 27304 39636
rect 30472 39627 30524 39636
rect 30472 39593 30481 39627
rect 30481 39593 30515 39627
rect 30515 39593 30524 39627
rect 30472 39584 30524 39593
rect 32680 39627 32732 39636
rect 32680 39593 32689 39627
rect 32689 39593 32723 39627
rect 32723 39593 32732 39627
rect 32680 39584 32732 39593
rect 34244 39584 34296 39636
rect 35440 39584 35492 39636
rect 39948 39584 40000 39636
rect 46572 39584 46624 39636
rect 48136 39627 48188 39636
rect 48136 39593 48145 39627
rect 48145 39593 48179 39627
rect 48179 39593 48188 39627
rect 48136 39584 48188 39593
rect 1400 39491 1452 39500
rect 1400 39457 1409 39491
rect 1409 39457 1443 39491
rect 1443 39457 1452 39491
rect 1400 39448 1452 39457
rect 2780 39491 2832 39500
rect 2780 39457 2789 39491
rect 2789 39457 2823 39491
rect 2823 39457 2832 39491
rect 2780 39448 2832 39457
rect 21272 39448 21324 39500
rect 22468 39491 22520 39500
rect 22468 39457 22477 39491
rect 22477 39457 22511 39491
rect 22511 39457 22520 39491
rect 22468 39448 22520 39457
rect 29828 39516 29880 39568
rect 37648 39516 37700 39568
rect 30564 39448 30616 39500
rect 26792 39380 26844 39432
rect 27252 39423 27304 39432
rect 27252 39389 27261 39423
rect 27261 39389 27295 39423
rect 27295 39389 27304 39423
rect 27252 39380 27304 39389
rect 28172 39423 28224 39432
rect 28172 39389 28181 39423
rect 28181 39389 28215 39423
rect 28215 39389 28224 39423
rect 28172 39380 28224 39389
rect 28264 39423 28316 39432
rect 28264 39389 28273 39423
rect 28273 39389 28307 39423
rect 28307 39389 28316 39423
rect 28264 39380 28316 39389
rect 31024 39380 31076 39432
rect 31392 39380 31444 39432
rect 1860 39312 1912 39364
rect 19432 39244 19484 39296
rect 20720 39312 20772 39364
rect 22560 39312 22612 39364
rect 25872 39312 25924 39364
rect 33600 39312 33652 39364
rect 35440 39380 35492 39432
rect 37832 39380 37884 39432
rect 38476 39380 38528 39432
rect 38844 39448 38896 39500
rect 40040 39448 40092 39500
rect 45376 39516 45428 39568
rect 42892 39491 42944 39500
rect 42892 39457 42901 39491
rect 42901 39457 42935 39491
rect 42935 39457 42944 39491
rect 42892 39448 42944 39457
rect 38752 39423 38804 39432
rect 38752 39389 38761 39423
rect 38761 39389 38795 39423
rect 38795 39389 38804 39423
rect 38752 39380 38804 39389
rect 39488 39380 39540 39432
rect 39856 39380 39908 39432
rect 40868 39380 40920 39432
rect 41052 39423 41104 39432
rect 41052 39389 41061 39423
rect 41061 39389 41095 39423
rect 41095 39389 41104 39423
rect 41052 39380 41104 39389
rect 42616 39423 42668 39432
rect 35256 39312 35308 39364
rect 23756 39244 23808 39296
rect 27068 39244 27120 39296
rect 27896 39244 27948 39296
rect 35348 39287 35400 39296
rect 35348 39253 35373 39287
rect 35373 39253 35400 39287
rect 35348 39244 35400 39253
rect 36728 39244 36780 39296
rect 38200 39244 38252 39296
rect 42340 39312 42392 39364
rect 40684 39244 40736 39296
rect 42616 39389 42625 39423
rect 42625 39389 42659 39423
rect 42659 39389 42668 39423
rect 42616 39380 42668 39389
rect 42800 39423 42852 39432
rect 42800 39389 42809 39423
rect 42809 39389 42843 39423
rect 42843 39389 42852 39423
rect 42800 39380 42852 39389
rect 43812 39380 43864 39432
rect 45100 39380 45152 39432
rect 46664 39448 46716 39500
rect 45652 39423 45704 39432
rect 45652 39389 45661 39423
rect 45661 39389 45695 39423
rect 45695 39389 45704 39423
rect 45652 39380 45704 39389
rect 46112 39423 46164 39432
rect 46112 39389 46121 39423
rect 46121 39389 46155 39423
rect 46155 39389 46164 39423
rect 46112 39380 46164 39389
rect 46848 39380 46900 39432
rect 48780 39423 48832 39432
rect 48780 39389 48789 39423
rect 48789 39389 48823 39423
rect 48823 39389 48832 39423
rect 48780 39380 48832 39389
rect 42524 39312 42576 39364
rect 43260 39244 43312 39296
rect 43444 39287 43496 39296
rect 43444 39253 43453 39287
rect 43453 39253 43487 39287
rect 43487 39253 43496 39287
rect 43444 39244 43496 39253
rect 44916 39244 44968 39296
rect 46020 39244 46072 39296
rect 48964 39244 49016 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 1860 39083 1912 39092
rect 1860 39049 1869 39083
rect 1869 39049 1903 39083
rect 1903 39049 1912 39083
rect 1860 39040 1912 39049
rect 19432 39040 19484 39092
rect 22560 39083 22612 39092
rect 22560 39049 22569 39083
rect 22569 39049 22603 39083
rect 22603 39049 22612 39083
rect 22560 39040 22612 39049
rect 3148 38904 3200 38956
rect 19984 38904 20036 38956
rect 20904 38947 20956 38956
rect 20904 38913 20913 38947
rect 20913 38913 20947 38947
rect 20947 38913 20956 38947
rect 20904 38904 20956 38913
rect 21088 38947 21140 38956
rect 21088 38913 21097 38947
rect 21097 38913 21131 38947
rect 21131 38913 21140 38947
rect 21088 38904 21140 38913
rect 23112 39040 23164 39092
rect 26240 39040 26292 39092
rect 27344 39040 27396 39092
rect 28172 39040 28224 39092
rect 31024 39083 31076 39092
rect 25228 38972 25280 39024
rect 31024 39049 31033 39083
rect 31033 39049 31067 39083
rect 31067 39049 31076 39083
rect 31024 39040 31076 39049
rect 35256 39083 35308 39092
rect 35256 39049 35265 39083
rect 35265 39049 35299 39083
rect 35299 39049 35308 39083
rect 35256 39040 35308 39049
rect 38476 39040 38528 39092
rect 40500 39083 40552 39092
rect 40500 39049 40509 39083
rect 40509 39049 40543 39083
rect 40543 39049 40552 39083
rect 40500 39040 40552 39049
rect 42524 39040 42576 39092
rect 43812 39083 43864 39092
rect 43812 39049 43821 39083
rect 43821 39049 43855 39083
rect 43855 39049 43864 39083
rect 43812 39040 43864 39049
rect 45100 39040 45152 39092
rect 45836 39040 45888 39092
rect 22744 38836 22796 38888
rect 23020 38947 23072 38956
rect 23020 38913 23029 38947
rect 23029 38913 23063 38947
rect 23063 38913 23072 38947
rect 23020 38904 23072 38913
rect 23112 38836 23164 38888
rect 23756 38904 23808 38956
rect 26240 38947 26292 38956
rect 26240 38913 26249 38947
rect 26249 38913 26283 38947
rect 26283 38913 26292 38947
rect 26240 38904 26292 38913
rect 27068 38947 27120 38956
rect 27068 38913 27077 38947
rect 27077 38913 27111 38947
rect 27111 38913 27120 38947
rect 27068 38904 27120 38913
rect 27712 38904 27764 38956
rect 24032 38879 24084 38888
rect 24032 38845 24041 38879
rect 24041 38845 24075 38879
rect 24075 38845 24084 38879
rect 24032 38836 24084 38845
rect 25596 38879 25648 38888
rect 25596 38845 25605 38879
rect 25605 38845 25639 38879
rect 25639 38845 25648 38879
rect 25596 38836 25648 38845
rect 30840 38904 30892 38956
rect 32312 38947 32364 38956
rect 32312 38913 32321 38947
rect 32321 38913 32355 38947
rect 32355 38913 32364 38947
rect 32312 38904 32364 38913
rect 33416 38947 33468 38956
rect 33416 38913 33425 38947
rect 33425 38913 33459 38947
rect 33459 38913 33468 38947
rect 33416 38904 33468 38913
rect 35808 38947 35860 38956
rect 33600 38879 33652 38888
rect 33600 38845 33609 38879
rect 33609 38845 33643 38879
rect 33643 38845 33652 38879
rect 33600 38836 33652 38845
rect 35808 38913 35817 38947
rect 35817 38913 35851 38947
rect 35851 38913 35860 38947
rect 35808 38904 35860 38913
rect 36728 38947 36780 38956
rect 36728 38913 36737 38947
rect 36737 38913 36771 38947
rect 36771 38913 36780 38947
rect 36728 38904 36780 38913
rect 39856 38972 39908 39024
rect 41052 38972 41104 39024
rect 43260 38972 43312 39024
rect 38200 38947 38252 38956
rect 38200 38913 38234 38947
rect 38234 38913 38252 38947
rect 38200 38904 38252 38913
rect 40684 38947 40736 38956
rect 40684 38913 40693 38947
rect 40693 38913 40727 38947
rect 40727 38913 40736 38947
rect 40684 38904 40736 38913
rect 41420 38947 41472 38956
rect 41420 38913 41429 38947
rect 41429 38913 41463 38947
rect 41463 38913 41472 38947
rect 41420 38904 41472 38913
rect 42340 38904 42392 38956
rect 42892 38947 42944 38956
rect 42892 38913 42901 38947
rect 42901 38913 42935 38947
rect 42935 38913 42944 38947
rect 42892 38904 42944 38913
rect 43352 38904 43404 38956
rect 43720 38972 43772 39024
rect 45192 38972 45244 39024
rect 46664 38972 46716 39024
rect 48964 39015 49016 39024
rect 48964 38981 48973 39015
rect 48973 38981 49007 39015
rect 49007 38981 49016 39015
rect 48964 38972 49016 38981
rect 44916 38947 44968 38956
rect 44916 38913 44950 38947
rect 44950 38913 44968 38947
rect 34428 38879 34480 38888
rect 34428 38845 34462 38879
rect 34462 38845 34480 38879
rect 34428 38836 34480 38845
rect 34796 38836 34848 38888
rect 35348 38836 35400 38888
rect 42800 38879 42852 38888
rect 42800 38845 42809 38879
rect 42809 38845 42843 38879
rect 42843 38845 42852 38879
rect 42800 38836 42852 38845
rect 33876 38768 33928 38820
rect 34060 38811 34112 38820
rect 34060 38777 34069 38811
rect 34069 38777 34103 38811
rect 34103 38777 34112 38811
rect 34060 38768 34112 38777
rect 42708 38768 42760 38820
rect 44916 38904 44968 38913
rect 48044 38904 48096 38956
rect 44088 38836 44140 38888
rect 50620 38879 50672 38888
rect 50620 38845 50629 38879
rect 50629 38845 50663 38879
rect 50663 38845 50672 38879
rect 50620 38836 50672 38845
rect 21180 38700 21232 38752
rect 32312 38700 32364 38752
rect 32864 38700 32916 38752
rect 34428 38700 34480 38752
rect 35992 38743 36044 38752
rect 35992 38709 36001 38743
rect 36001 38709 36035 38743
rect 36035 38709 36044 38743
rect 35992 38700 36044 38709
rect 36544 38743 36596 38752
rect 36544 38709 36553 38743
rect 36553 38709 36587 38743
rect 36587 38709 36596 38743
rect 36544 38700 36596 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 65654 38598 65706 38650
rect 65718 38598 65770 38650
rect 65782 38598 65834 38650
rect 65846 38598 65898 38650
rect 65910 38598 65962 38650
rect 3240 38496 3292 38548
rect 20720 38496 20772 38548
rect 24032 38496 24084 38548
rect 27712 38539 27764 38548
rect 27712 38505 27721 38539
rect 27721 38505 27755 38539
rect 27755 38505 27764 38539
rect 27712 38496 27764 38505
rect 32864 38496 32916 38548
rect 35440 38496 35492 38548
rect 39856 38496 39908 38548
rect 45192 38496 45244 38548
rect 44088 38428 44140 38480
rect 37372 38403 37424 38412
rect 37372 38369 37381 38403
rect 37381 38369 37415 38403
rect 37415 38369 37424 38403
rect 37372 38360 37424 38369
rect 45836 38403 45888 38412
rect 45836 38369 45845 38403
rect 45845 38369 45879 38403
rect 45879 38369 45888 38403
rect 45836 38360 45888 38369
rect 46020 38403 46072 38412
rect 46020 38369 46029 38403
rect 46029 38369 46063 38403
rect 46063 38369 46072 38403
rect 46020 38360 46072 38369
rect 19984 38292 20036 38344
rect 22376 38292 22428 38344
rect 23388 38292 23440 38344
rect 24400 38335 24452 38344
rect 24400 38301 24409 38335
rect 24409 38301 24443 38335
rect 24443 38301 24452 38335
rect 24400 38292 24452 38301
rect 27896 38335 27948 38344
rect 27896 38301 27905 38335
rect 27905 38301 27939 38335
rect 27939 38301 27948 38335
rect 27896 38292 27948 38301
rect 30196 38292 30248 38344
rect 30840 38335 30892 38344
rect 30840 38301 30849 38335
rect 30849 38301 30883 38335
rect 30883 38301 30892 38335
rect 30840 38292 30892 38301
rect 21180 38267 21232 38276
rect 21180 38233 21214 38267
rect 21214 38233 21232 38267
rect 21180 38224 21232 38233
rect 24676 38267 24728 38276
rect 24676 38233 24710 38267
rect 24710 38233 24728 38267
rect 24676 38224 24728 38233
rect 32128 38224 32180 38276
rect 33784 38267 33836 38276
rect 33784 38233 33793 38267
rect 33793 38233 33827 38267
rect 33827 38233 33836 38267
rect 33784 38224 33836 38233
rect 34060 38224 34112 38276
rect 34520 38224 34572 38276
rect 36544 38292 36596 38344
rect 37648 38335 37700 38344
rect 37648 38301 37657 38335
rect 37657 38301 37691 38335
rect 37691 38301 37700 38335
rect 37648 38292 37700 38301
rect 38384 38292 38436 38344
rect 40960 38292 41012 38344
rect 43444 38292 43496 38344
rect 35992 38224 36044 38276
rect 40592 38267 40644 38276
rect 40592 38233 40601 38267
rect 40601 38233 40635 38267
rect 40635 38233 40644 38267
rect 40592 38224 40644 38233
rect 66812 38292 66864 38344
rect 19984 38156 20036 38208
rect 20904 38156 20956 38208
rect 27252 38156 27304 38208
rect 29644 38199 29696 38208
rect 29644 38165 29653 38199
rect 29653 38165 29687 38199
rect 29687 38165 29696 38199
rect 29644 38156 29696 38165
rect 32220 38156 32272 38208
rect 47584 38224 47636 38276
rect 50068 38156 50120 38208
rect 66628 38156 66680 38208
rect 66812 38156 66864 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 20904 37952 20956 38004
rect 24400 37952 24452 38004
rect 32128 37995 32180 38004
rect 32128 37961 32137 37995
rect 32137 37961 32171 37995
rect 32171 37961 32180 37995
rect 32128 37952 32180 37961
rect 38568 37952 38620 38004
rect 40868 37952 40920 38004
rect 19984 37884 20036 37936
rect 27160 37927 27212 37936
rect 27160 37893 27169 37927
rect 27169 37893 27203 37927
rect 27203 37893 27212 37927
rect 27160 37884 27212 37893
rect 28816 37884 28868 37936
rect 29644 37927 29696 37936
rect 29644 37893 29678 37927
rect 29678 37893 29696 37927
rect 29644 37884 29696 37893
rect 37464 37884 37516 37936
rect 38752 37927 38804 37936
rect 38752 37893 38761 37927
rect 38761 37893 38795 37927
rect 38795 37893 38804 37927
rect 38752 37884 38804 37893
rect 39948 37884 40000 37936
rect 23296 37859 23348 37868
rect 23296 37825 23305 37859
rect 23305 37825 23339 37859
rect 23339 37825 23348 37859
rect 23296 37816 23348 37825
rect 25780 37816 25832 37868
rect 26056 37859 26108 37868
rect 26056 37825 26065 37859
rect 26065 37825 26099 37859
rect 26099 37825 26108 37859
rect 26056 37816 26108 37825
rect 26424 37816 26476 37868
rect 29368 37859 29420 37868
rect 29368 37825 29377 37859
rect 29377 37825 29411 37859
rect 29411 37825 29420 37859
rect 29368 37816 29420 37825
rect 32312 37859 32364 37868
rect 32312 37825 32321 37859
rect 32321 37825 32355 37859
rect 32355 37825 32364 37859
rect 32312 37816 32364 37825
rect 32680 37816 32732 37868
rect 33324 37816 33376 37868
rect 35808 37816 35860 37868
rect 37556 37859 37608 37868
rect 37556 37825 37565 37859
rect 37565 37825 37599 37859
rect 37599 37825 37608 37859
rect 37556 37816 37608 37825
rect 39008 37859 39060 37868
rect 39008 37825 39017 37859
rect 39017 37825 39051 37859
rect 39051 37825 39060 37859
rect 39008 37816 39060 37825
rect 24216 37791 24268 37800
rect 20 37680 72 37732
rect 24216 37757 24225 37791
rect 24225 37757 24259 37791
rect 24259 37757 24268 37791
rect 24216 37748 24268 37757
rect 26148 37748 26200 37800
rect 33232 37748 33284 37800
rect 34704 37748 34756 37800
rect 39488 37816 39540 37868
rect 39856 37859 39908 37868
rect 39856 37825 39865 37859
rect 39865 37825 39899 37859
rect 39899 37825 39908 37859
rect 39856 37816 39908 37825
rect 44364 37927 44416 37936
rect 44364 37893 44373 37927
rect 44373 37893 44407 37927
rect 44407 37893 44416 37927
rect 44364 37884 44416 37893
rect 47308 37884 47360 37936
rect 48044 37884 48096 37936
rect 50068 37927 50120 37936
rect 50068 37893 50077 37927
rect 50077 37893 50111 37927
rect 50111 37893 50120 37927
rect 50068 37884 50120 37893
rect 42708 37859 42760 37868
rect 42708 37825 42717 37859
rect 42717 37825 42751 37859
rect 42751 37825 42760 37859
rect 42708 37816 42760 37825
rect 45008 37859 45060 37868
rect 45008 37825 45017 37859
rect 45017 37825 45051 37859
rect 45051 37825 45060 37859
rect 45008 37816 45060 37825
rect 25320 37612 25372 37664
rect 27344 37655 27396 37664
rect 27344 37621 27353 37655
rect 27353 37621 27387 37655
rect 27387 37621 27396 37655
rect 27344 37612 27396 37621
rect 27528 37655 27580 37664
rect 27528 37621 27537 37655
rect 27537 37621 27571 37655
rect 27571 37621 27580 37655
rect 27528 37612 27580 37621
rect 30012 37612 30064 37664
rect 35440 37680 35492 37732
rect 39028 37680 39080 37732
rect 39304 37748 39356 37800
rect 46572 37748 46624 37800
rect 47768 37791 47820 37800
rect 47768 37757 47777 37791
rect 47777 37757 47811 37791
rect 47811 37757 47820 37791
rect 47768 37748 47820 37757
rect 48044 37791 48096 37800
rect 48044 37757 48053 37791
rect 48053 37757 48087 37791
rect 48087 37757 48096 37791
rect 48044 37748 48096 37757
rect 51724 37791 51776 37800
rect 39856 37680 39908 37732
rect 51724 37757 51733 37791
rect 51733 37757 51767 37791
rect 51767 37757 51776 37791
rect 51724 37748 51776 37757
rect 30380 37612 30432 37664
rect 38936 37612 38988 37664
rect 44916 37612 44968 37664
rect 46848 37612 46900 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 27252 37408 27304 37460
rect 37556 37408 37608 37460
rect 39304 37408 39356 37460
rect 39488 37408 39540 37460
rect 40684 37408 40736 37460
rect 47768 37408 47820 37460
rect 3240 37136 3292 37188
rect 25320 37315 25372 37324
rect 25320 37281 25329 37315
rect 25329 37281 25363 37315
rect 25363 37281 25372 37315
rect 25320 37272 25372 37281
rect 27712 37340 27764 37392
rect 27896 37340 27948 37392
rect 30012 37340 30064 37392
rect 27160 37315 27212 37324
rect 27160 37281 27169 37315
rect 27169 37281 27203 37315
rect 27203 37281 27212 37315
rect 27160 37272 27212 37281
rect 27252 37272 27304 37324
rect 35440 37315 35492 37324
rect 35440 37281 35449 37315
rect 35449 37281 35483 37315
rect 35483 37281 35492 37315
rect 35440 37272 35492 37281
rect 35624 37272 35676 37324
rect 35992 37272 36044 37324
rect 39120 37315 39172 37324
rect 22744 37136 22796 37188
rect 26608 37136 26660 37188
rect 22928 37068 22980 37120
rect 24860 37111 24912 37120
rect 24860 37077 24869 37111
rect 24869 37077 24903 37111
rect 24903 37077 24912 37111
rect 24860 37068 24912 37077
rect 25504 37068 25556 37120
rect 28080 37247 28132 37256
rect 28080 37213 28089 37247
rect 28089 37213 28123 37247
rect 28123 37213 28132 37247
rect 28356 37247 28408 37256
rect 28080 37204 28132 37213
rect 28356 37213 28365 37247
rect 28365 37213 28399 37247
rect 28399 37213 28408 37247
rect 28356 37204 28408 37213
rect 30012 37247 30064 37256
rect 30012 37213 30021 37247
rect 30021 37213 30055 37247
rect 30055 37213 30064 37247
rect 30012 37204 30064 37213
rect 32772 37247 32824 37256
rect 32772 37213 32781 37247
rect 32781 37213 32815 37247
rect 32815 37213 32824 37247
rect 32772 37204 32824 37213
rect 33508 37204 33560 37256
rect 35808 37204 35860 37256
rect 39120 37281 39129 37315
rect 39129 37281 39163 37315
rect 39163 37281 39172 37315
rect 39120 37272 39172 37281
rect 39580 37272 39632 37324
rect 38936 37247 38988 37256
rect 38936 37213 38945 37247
rect 38945 37213 38979 37247
rect 38979 37213 38988 37247
rect 38936 37204 38988 37213
rect 39028 37247 39080 37256
rect 39028 37213 39037 37247
rect 39037 37213 39071 37247
rect 39071 37213 39080 37247
rect 39028 37204 39080 37213
rect 39396 37204 39448 37256
rect 39488 37204 39540 37256
rect 40868 37204 40920 37256
rect 43076 37340 43128 37392
rect 41880 37247 41932 37256
rect 41880 37213 41889 37247
rect 41889 37213 41923 37247
rect 41923 37213 41932 37247
rect 41880 37204 41932 37213
rect 42800 37204 42852 37256
rect 44364 37204 44416 37256
rect 45192 37247 45244 37256
rect 45192 37213 45201 37247
rect 45201 37213 45235 37247
rect 45235 37213 45244 37247
rect 45192 37204 45244 37213
rect 46848 37204 46900 37256
rect 29828 37068 29880 37120
rect 30380 37068 30432 37120
rect 33876 37068 33928 37120
rect 43260 37136 43312 37188
rect 44732 37136 44784 37188
rect 44824 37136 44876 37188
rect 35992 37068 36044 37120
rect 45008 37068 45060 37120
rect 46572 37111 46624 37120
rect 46572 37077 46581 37111
rect 46581 37077 46615 37111
rect 46615 37077 46624 37111
rect 46572 37068 46624 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 22744 36907 22796 36916
rect 22744 36873 22753 36907
rect 22753 36873 22787 36907
rect 22787 36873 22796 36907
rect 22744 36864 22796 36873
rect 24676 36907 24728 36916
rect 24676 36873 24685 36907
rect 24685 36873 24719 36907
rect 24719 36873 24728 36907
rect 24676 36864 24728 36873
rect 29736 36864 29788 36916
rect 30012 36907 30064 36916
rect 30012 36873 30037 36907
rect 30037 36873 30064 36907
rect 30196 36907 30248 36916
rect 30012 36864 30064 36873
rect 30196 36873 30205 36907
rect 30205 36873 30239 36907
rect 30239 36873 30248 36907
rect 30196 36864 30248 36873
rect 25688 36796 25740 36848
rect 29828 36839 29880 36848
rect 29828 36805 29837 36839
rect 29837 36805 29871 36839
rect 29871 36805 29880 36839
rect 29828 36796 29880 36805
rect 23296 36728 23348 36780
rect 24860 36771 24912 36780
rect 24860 36737 24869 36771
rect 24869 36737 24903 36771
rect 24903 36737 24912 36771
rect 24860 36728 24912 36737
rect 25504 36728 25556 36780
rect 32680 36796 32732 36848
rect 30196 36728 30248 36780
rect 1584 36524 1636 36576
rect 26240 36660 26292 36712
rect 24308 36524 24360 36576
rect 27344 36660 27396 36712
rect 28816 36703 28868 36712
rect 28816 36669 28825 36703
rect 28825 36669 28859 36703
rect 28859 36669 28868 36703
rect 28816 36660 28868 36669
rect 31392 36660 31444 36712
rect 29552 36592 29604 36644
rect 33324 36728 33376 36780
rect 33876 36771 33928 36780
rect 33876 36737 33885 36771
rect 33885 36737 33919 36771
rect 33919 36737 33928 36771
rect 33876 36728 33928 36737
rect 36176 36839 36228 36848
rect 36176 36805 36185 36839
rect 36185 36805 36219 36839
rect 36219 36805 36228 36839
rect 36176 36796 36228 36805
rect 37832 36864 37884 36916
rect 38384 36864 38436 36916
rect 38936 36864 38988 36916
rect 35808 36728 35860 36780
rect 40592 36796 40644 36848
rect 37372 36771 37424 36780
rect 37372 36737 37381 36771
rect 37381 36737 37415 36771
rect 37415 36737 37424 36771
rect 37372 36728 37424 36737
rect 38384 36771 38436 36780
rect 34796 36703 34848 36712
rect 34796 36669 34805 36703
rect 34805 36669 34839 36703
rect 34839 36669 34848 36703
rect 34796 36660 34848 36669
rect 34888 36703 34940 36712
rect 34888 36669 34922 36703
rect 34922 36669 34940 36703
rect 34888 36660 34940 36669
rect 35440 36660 35492 36712
rect 38384 36737 38393 36771
rect 38393 36737 38427 36771
rect 38427 36737 38436 36771
rect 38384 36728 38436 36737
rect 39028 36771 39080 36780
rect 39028 36737 39037 36771
rect 39037 36737 39071 36771
rect 39071 36737 39080 36771
rect 39028 36728 39080 36737
rect 39212 36771 39264 36780
rect 39212 36737 39221 36771
rect 39221 36737 39255 36771
rect 39255 36737 39264 36771
rect 39212 36728 39264 36737
rect 41880 36728 41932 36780
rect 42708 36864 42760 36916
rect 43352 36864 43404 36916
rect 44824 36907 44876 36916
rect 44824 36873 44833 36907
rect 44833 36873 44867 36907
rect 44867 36873 44876 36907
rect 44824 36864 44876 36873
rect 44916 36864 44968 36916
rect 45376 36864 45428 36916
rect 42432 36796 42484 36848
rect 43260 36771 43312 36780
rect 43260 36737 43269 36771
rect 43269 36737 43303 36771
rect 43303 36737 43312 36771
rect 43260 36728 43312 36737
rect 44824 36728 44876 36780
rect 34520 36635 34572 36644
rect 34520 36601 34529 36635
rect 34529 36601 34563 36635
rect 34563 36601 34572 36635
rect 34520 36592 34572 36601
rect 42708 36660 42760 36712
rect 43352 36703 43404 36712
rect 42800 36592 42852 36644
rect 43352 36669 43361 36703
rect 43361 36669 43395 36703
rect 43395 36669 43404 36703
rect 43352 36660 43404 36669
rect 44916 36660 44968 36712
rect 44732 36592 44784 36644
rect 45192 36592 45244 36644
rect 29920 36524 29972 36576
rect 30472 36524 30524 36576
rect 35532 36524 35584 36576
rect 35716 36524 35768 36576
rect 36544 36567 36596 36576
rect 36544 36533 36553 36567
rect 36553 36533 36587 36567
rect 36587 36533 36596 36567
rect 36544 36524 36596 36533
rect 40408 36524 40460 36576
rect 41328 36567 41380 36576
rect 41328 36533 41337 36567
rect 41337 36533 41371 36567
rect 41371 36533 41380 36567
rect 41328 36524 41380 36533
rect 45652 36728 45704 36780
rect 46388 36771 46440 36780
rect 46388 36737 46397 36771
rect 46397 36737 46431 36771
rect 46431 36737 46440 36771
rect 46388 36728 46440 36737
rect 46756 36728 46808 36780
rect 47860 36660 47912 36712
rect 46756 36592 46808 36644
rect 46572 36524 46624 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 26608 36363 26660 36372
rect 26608 36329 26617 36363
rect 26617 36329 26651 36363
rect 26651 36329 26660 36363
rect 26608 36320 26660 36329
rect 32312 36363 32364 36372
rect 32312 36329 32321 36363
rect 32321 36329 32355 36363
rect 32355 36329 32364 36363
rect 32312 36320 32364 36329
rect 33232 36320 33284 36372
rect 33508 36363 33560 36372
rect 33508 36329 33517 36363
rect 33517 36329 33551 36363
rect 33551 36329 33560 36363
rect 33508 36320 33560 36329
rect 36176 36320 36228 36372
rect 39212 36320 39264 36372
rect 41328 36320 41380 36372
rect 46388 36320 46440 36372
rect 47860 36363 47912 36372
rect 47860 36329 47869 36363
rect 47869 36329 47903 36363
rect 47903 36329 47912 36363
rect 47860 36320 47912 36329
rect 1584 36227 1636 36236
rect 1584 36193 1593 36227
rect 1593 36193 1627 36227
rect 1627 36193 1636 36227
rect 1584 36184 1636 36193
rect 2780 36227 2832 36236
rect 2780 36193 2789 36227
rect 2789 36193 2823 36227
rect 2823 36193 2832 36227
rect 2780 36184 2832 36193
rect 28080 36184 28132 36236
rect 1400 36159 1452 36168
rect 1400 36125 1409 36159
rect 1409 36125 1443 36159
rect 1443 36125 1452 36159
rect 1400 36116 1452 36125
rect 22284 36159 22336 36168
rect 22284 36125 22293 36159
rect 22293 36125 22327 36159
rect 22327 36125 22336 36159
rect 22284 36116 22336 36125
rect 23572 36116 23624 36168
rect 25780 36116 25832 36168
rect 27528 36116 27580 36168
rect 28448 36116 28500 36168
rect 23020 36048 23072 36100
rect 29920 36116 29972 36168
rect 30840 36184 30892 36236
rect 35992 36227 36044 36236
rect 35992 36193 36001 36227
rect 36001 36193 36035 36227
rect 36035 36193 36044 36227
rect 35992 36184 36044 36193
rect 39028 36184 39080 36236
rect 44824 36184 44876 36236
rect 34704 36116 34756 36168
rect 37924 36159 37976 36168
rect 37924 36125 37933 36159
rect 37933 36125 37967 36159
rect 37967 36125 37976 36159
rect 37924 36116 37976 36125
rect 39764 36116 39816 36168
rect 42432 36116 42484 36168
rect 42984 36116 43036 36168
rect 45560 36116 45612 36168
rect 46572 36116 46624 36168
rect 66904 36116 66956 36168
rect 31300 36048 31352 36100
rect 33876 36048 33928 36100
rect 36360 36048 36412 36100
rect 38936 36048 38988 36100
rect 23756 35980 23808 36032
rect 25320 36023 25372 36032
rect 25320 35989 25329 36023
rect 25329 35989 25363 36023
rect 25363 35989 25372 36023
rect 25320 35980 25372 35989
rect 28724 36023 28776 36032
rect 28724 35989 28733 36023
rect 28733 35989 28767 36023
rect 28767 35989 28776 36023
rect 28724 35980 28776 35989
rect 29552 36023 29604 36032
rect 29552 35989 29561 36023
rect 29561 35989 29595 36023
rect 29595 35989 29604 36023
rect 29552 35980 29604 35989
rect 33324 36023 33376 36032
rect 33324 35989 33349 36023
rect 33349 35989 33376 36023
rect 33324 35980 33376 35989
rect 44180 35980 44232 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 14464 35708 14516 35760
rect 1400 35640 1452 35692
rect 19156 35683 19208 35692
rect 19156 35649 19165 35683
rect 19165 35649 19199 35683
rect 19199 35649 19208 35683
rect 19156 35640 19208 35649
rect 19984 35640 20036 35692
rect 20720 35683 20772 35692
rect 20720 35649 20729 35683
rect 20729 35649 20763 35683
rect 20763 35649 20772 35683
rect 20720 35640 20772 35649
rect 22652 35683 22704 35692
rect 8024 35504 8076 35556
rect 20352 35572 20404 35624
rect 20904 35615 20956 35624
rect 20904 35581 20913 35615
rect 20913 35581 20947 35615
rect 20947 35581 20956 35615
rect 20904 35572 20956 35581
rect 1676 35436 1728 35488
rect 14464 35436 14516 35488
rect 22652 35649 22661 35683
rect 22661 35649 22695 35683
rect 22695 35649 22704 35683
rect 22652 35640 22704 35649
rect 36176 35776 36228 35828
rect 36360 35819 36412 35828
rect 36360 35785 36369 35819
rect 36369 35785 36403 35819
rect 36403 35785 36412 35819
rect 36360 35776 36412 35785
rect 37924 35776 37976 35828
rect 25320 35708 25372 35760
rect 29552 35708 29604 35760
rect 24492 35683 24544 35692
rect 24492 35649 24526 35683
rect 24526 35649 24544 35683
rect 24492 35640 24544 35649
rect 27436 35640 27488 35692
rect 28724 35640 28776 35692
rect 30748 35640 30800 35692
rect 32312 35708 32364 35760
rect 67364 35776 67416 35828
rect 42432 35751 42484 35760
rect 31392 35683 31444 35692
rect 31392 35649 31401 35683
rect 31401 35649 31435 35683
rect 31435 35649 31444 35683
rect 32404 35683 32456 35692
rect 31392 35640 31444 35649
rect 22560 35572 22612 35624
rect 32404 35649 32413 35683
rect 32413 35649 32447 35683
rect 32447 35649 32456 35683
rect 32404 35640 32456 35649
rect 33416 35640 33468 35692
rect 25688 35436 25740 35488
rect 26976 35479 27028 35488
rect 26976 35445 26985 35479
rect 26985 35445 27019 35479
rect 27019 35445 27028 35479
rect 26976 35436 27028 35445
rect 30012 35479 30064 35488
rect 30012 35445 30021 35479
rect 30021 35445 30055 35479
rect 30055 35445 30064 35479
rect 30012 35436 30064 35445
rect 42432 35717 42441 35751
rect 42441 35717 42475 35751
rect 42475 35717 42484 35751
rect 42432 35708 42484 35717
rect 42800 35751 42852 35760
rect 42800 35717 42809 35751
rect 42809 35717 42843 35751
rect 42843 35717 42852 35751
rect 42800 35708 42852 35717
rect 35624 35683 35676 35692
rect 35624 35649 35633 35683
rect 35633 35649 35667 35683
rect 35667 35649 35676 35683
rect 35624 35640 35676 35649
rect 36544 35683 36596 35692
rect 36544 35649 36553 35683
rect 36553 35649 36587 35683
rect 36587 35649 36596 35683
rect 36544 35640 36596 35649
rect 37280 35640 37332 35692
rect 38016 35640 38068 35692
rect 39212 35683 39264 35692
rect 39212 35649 39221 35683
rect 39221 35649 39255 35683
rect 39255 35649 39264 35683
rect 39212 35640 39264 35649
rect 40316 35640 40368 35692
rect 41604 35640 41656 35692
rect 35992 35572 36044 35624
rect 40500 35615 40552 35624
rect 40500 35581 40509 35615
rect 40509 35581 40543 35615
rect 40543 35581 40552 35615
rect 40500 35572 40552 35581
rect 43996 35640 44048 35692
rect 46848 35683 46900 35692
rect 46848 35649 46857 35683
rect 46857 35649 46891 35683
rect 46891 35649 46900 35683
rect 46848 35640 46900 35649
rect 47860 35640 47912 35692
rect 66904 35708 66956 35760
rect 35348 35504 35400 35556
rect 42800 35572 42852 35624
rect 43444 35615 43496 35624
rect 43444 35581 43453 35615
rect 43453 35581 43487 35615
rect 43487 35581 43496 35615
rect 43444 35572 43496 35581
rect 49608 35615 49660 35624
rect 49608 35581 49617 35615
rect 49617 35581 49651 35615
rect 49651 35581 49660 35615
rect 49608 35572 49660 35581
rect 65984 35615 66036 35624
rect 65984 35581 65993 35615
rect 65993 35581 66027 35615
rect 66027 35581 66036 35615
rect 65984 35572 66036 35581
rect 67548 35615 67600 35624
rect 67548 35581 67557 35615
rect 67557 35581 67591 35615
rect 67591 35581 67600 35615
rect 67548 35572 67600 35581
rect 44824 35547 44876 35556
rect 44824 35513 44833 35547
rect 44833 35513 44867 35547
rect 44867 35513 44876 35547
rect 44824 35504 44876 35513
rect 31484 35436 31536 35488
rect 32588 35479 32640 35488
rect 32588 35445 32597 35479
rect 32597 35445 32631 35479
rect 32631 35445 32640 35479
rect 32588 35436 32640 35445
rect 33140 35479 33192 35488
rect 33140 35445 33149 35479
rect 33149 35445 33183 35479
rect 33183 35445 33192 35479
rect 33140 35436 33192 35445
rect 35440 35436 35492 35488
rect 35532 35436 35584 35488
rect 35900 35436 35952 35488
rect 39120 35436 39172 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 20076 35232 20128 35284
rect 21732 35232 21784 35284
rect 22284 35275 22336 35284
rect 22284 35241 22293 35275
rect 22293 35241 22327 35275
rect 22327 35241 22336 35275
rect 22284 35232 22336 35241
rect 23020 35275 23072 35284
rect 23020 35241 23029 35275
rect 23029 35241 23063 35275
rect 23063 35241 23072 35275
rect 23020 35232 23072 35241
rect 22652 35164 22704 35216
rect 25688 35232 25740 35284
rect 27068 35096 27120 35148
rect 27712 35164 27764 35216
rect 29920 35275 29972 35284
rect 29920 35241 29929 35275
rect 29929 35241 29963 35275
rect 29963 35241 29972 35275
rect 29920 35232 29972 35241
rect 31300 35275 31352 35284
rect 31300 35241 31309 35275
rect 31309 35241 31343 35275
rect 31343 35241 31352 35275
rect 31300 35232 31352 35241
rect 31576 35232 31628 35284
rect 30472 35164 30524 35216
rect 34520 35164 34572 35216
rect 32588 35139 32640 35148
rect 20812 35071 20864 35080
rect 20812 35037 20821 35071
rect 20821 35037 20855 35071
rect 20855 35037 20864 35071
rect 20812 35028 20864 35037
rect 22376 35071 22428 35080
rect 22376 35037 22385 35071
rect 22385 35037 22419 35071
rect 22419 35037 22428 35071
rect 22376 35028 22428 35037
rect 23756 35028 23808 35080
rect 25320 35071 25372 35080
rect 20536 35003 20588 35012
rect 20536 34969 20545 35003
rect 20545 34969 20579 35003
rect 20579 34969 20588 35003
rect 20536 34960 20588 34969
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 26976 35028 27028 35080
rect 25504 34960 25556 35012
rect 24860 34935 24912 34944
rect 24860 34901 24869 34935
rect 24869 34901 24903 34935
rect 24903 34901 24912 34935
rect 24860 34892 24912 34901
rect 32588 35105 32597 35139
rect 32597 35105 32631 35139
rect 32631 35105 32640 35139
rect 32588 35096 32640 35105
rect 35256 35096 35308 35148
rect 37372 35232 37424 35284
rect 38936 35275 38988 35284
rect 38936 35241 38945 35275
rect 38945 35241 38979 35275
rect 38979 35241 38988 35275
rect 38936 35232 38988 35241
rect 43444 35232 43496 35284
rect 65984 35232 66036 35284
rect 45652 35207 45704 35216
rect 35900 35139 35952 35148
rect 35900 35105 35909 35139
rect 35909 35105 35943 35139
rect 35943 35105 35952 35139
rect 35900 35096 35952 35105
rect 40132 35139 40184 35148
rect 40132 35105 40141 35139
rect 40141 35105 40175 35139
rect 40175 35105 40184 35139
rect 40132 35096 40184 35105
rect 40316 35096 40368 35148
rect 45652 35173 45661 35207
rect 45661 35173 45695 35207
rect 45695 35173 45704 35207
rect 45652 35164 45704 35173
rect 42800 35139 42852 35148
rect 42800 35105 42809 35139
rect 42809 35105 42843 35139
rect 42843 35105 42852 35139
rect 42800 35096 42852 35105
rect 49240 35139 49292 35148
rect 49240 35105 49249 35139
rect 49249 35105 49283 35139
rect 49283 35105 49292 35139
rect 49240 35096 49292 35105
rect 28080 35071 28132 35080
rect 28080 35037 28089 35071
rect 28089 35037 28123 35071
rect 28123 35037 28132 35071
rect 28356 35071 28408 35080
rect 28080 35028 28132 35037
rect 28356 35037 28365 35071
rect 28365 35037 28399 35071
rect 28399 35037 28408 35071
rect 28356 35028 28408 35037
rect 30012 34960 30064 35012
rect 30840 35028 30892 35080
rect 31484 35071 31536 35080
rect 31484 35037 31493 35071
rect 31493 35037 31527 35071
rect 31527 35037 31536 35071
rect 31484 35028 31536 35037
rect 33140 35028 33192 35080
rect 33968 35028 34020 35080
rect 35624 35071 35676 35080
rect 35624 35037 35633 35071
rect 35633 35037 35667 35071
rect 35667 35037 35676 35071
rect 35624 35028 35676 35037
rect 38936 35028 38988 35080
rect 39120 35071 39172 35080
rect 39120 35037 39129 35071
rect 39129 35037 39163 35071
rect 39163 35037 39172 35071
rect 39120 35028 39172 35037
rect 42984 35071 43036 35080
rect 42984 35037 42993 35071
rect 42993 35037 43027 35071
rect 43027 35037 43036 35071
rect 42984 35028 43036 35037
rect 29736 34935 29788 34944
rect 29736 34901 29761 34935
rect 29761 34901 29788 34935
rect 29736 34892 29788 34901
rect 30196 34892 30248 34944
rect 33968 34935 34020 34944
rect 33968 34901 33977 34935
rect 33977 34901 34011 34935
rect 34011 34901 34020 34935
rect 33968 34892 34020 34901
rect 37464 34960 37516 35012
rect 40960 34960 41012 35012
rect 44272 35028 44324 35080
rect 45284 35028 45336 35080
rect 47492 35071 47544 35080
rect 47492 35037 47501 35071
rect 47501 35037 47535 35071
rect 47535 35037 47544 35071
rect 47492 35028 47544 35037
rect 67456 35071 67508 35080
rect 67456 35037 67465 35071
rect 67465 35037 67499 35071
rect 67499 35037 67508 35071
rect 67456 35028 67508 35037
rect 47676 35003 47728 35012
rect 47676 34969 47685 35003
rect 47685 34969 47719 35003
rect 47719 34969 47728 35003
rect 47676 34960 47728 34969
rect 38016 34892 38068 34944
rect 38108 34892 38160 34944
rect 41788 34892 41840 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 24492 34688 24544 34740
rect 25320 34688 25372 34740
rect 27436 34731 27488 34740
rect 27436 34697 27445 34731
rect 27445 34697 27479 34731
rect 27479 34697 27488 34731
rect 27436 34688 27488 34697
rect 31576 34731 31628 34740
rect 31576 34697 31585 34731
rect 31585 34697 31619 34731
rect 31619 34697 31628 34731
rect 31576 34688 31628 34697
rect 27068 34663 27120 34672
rect 27068 34629 27077 34663
rect 27077 34629 27111 34663
rect 27111 34629 27120 34663
rect 27068 34620 27120 34629
rect 28816 34620 28868 34672
rect 33416 34731 33468 34740
rect 33416 34697 33425 34731
rect 33425 34697 33459 34731
rect 33459 34697 33468 34731
rect 33416 34688 33468 34697
rect 35256 34688 35308 34740
rect 40224 34688 40276 34740
rect 40500 34688 40552 34740
rect 41604 34731 41656 34740
rect 41604 34697 41613 34731
rect 41613 34697 41647 34731
rect 41647 34697 41656 34731
rect 41604 34688 41656 34697
rect 43996 34731 44048 34740
rect 43996 34697 44005 34731
rect 44005 34697 44039 34731
rect 44039 34697 44048 34731
rect 43996 34688 44048 34697
rect 45376 34688 45428 34740
rect 47492 34688 47544 34740
rect 47676 34731 47728 34740
rect 47676 34697 47685 34731
rect 47685 34697 47719 34731
rect 47719 34697 47728 34731
rect 47676 34688 47728 34697
rect 20536 34552 20588 34604
rect 23480 34552 23532 34604
rect 24860 34595 24912 34604
rect 24860 34561 24869 34595
rect 24869 34561 24903 34595
rect 24903 34561 24912 34595
rect 24860 34552 24912 34561
rect 26056 34552 26108 34604
rect 30196 34595 30248 34604
rect 30196 34561 30205 34595
rect 30205 34561 30239 34595
rect 30239 34561 30248 34595
rect 30196 34552 30248 34561
rect 32312 34595 32364 34604
rect 32312 34561 32321 34595
rect 32321 34561 32355 34595
rect 32355 34561 32364 34595
rect 32312 34552 32364 34561
rect 33232 34663 33284 34672
rect 33232 34629 33257 34663
rect 33257 34629 33284 34663
rect 37740 34663 37792 34672
rect 33232 34620 33284 34629
rect 37740 34629 37749 34663
rect 37749 34629 37783 34663
rect 37783 34629 37792 34663
rect 37740 34620 37792 34629
rect 33968 34552 34020 34604
rect 35348 34595 35400 34604
rect 35348 34561 35357 34595
rect 35357 34561 35391 34595
rect 35391 34561 35400 34595
rect 35348 34552 35400 34561
rect 35440 34552 35492 34604
rect 38016 34552 38068 34604
rect 39488 34552 39540 34604
rect 40960 34595 41012 34604
rect 40960 34561 40969 34595
rect 40969 34561 41003 34595
rect 41003 34561 41012 34595
rect 40960 34552 41012 34561
rect 41788 34595 41840 34604
rect 41788 34561 41797 34595
rect 41797 34561 41831 34595
rect 41831 34561 41840 34595
rect 41788 34552 41840 34561
rect 44180 34595 44232 34604
rect 44180 34561 44189 34595
rect 44189 34561 44223 34595
rect 44223 34561 44232 34595
rect 44180 34552 44232 34561
rect 45560 34552 45612 34604
rect 45744 34595 45796 34604
rect 45744 34561 45778 34595
rect 45778 34561 45796 34595
rect 45744 34552 45796 34561
rect 46756 34552 46808 34604
rect 67272 34595 67324 34604
rect 67272 34561 67281 34595
rect 67281 34561 67315 34595
rect 67315 34561 67324 34595
rect 67272 34552 67324 34561
rect 1400 34527 1452 34536
rect 1400 34493 1409 34527
rect 1409 34493 1443 34527
rect 1443 34493 1452 34527
rect 1400 34484 1452 34493
rect 39120 34527 39172 34536
rect 39120 34493 39129 34527
rect 39129 34493 39163 34527
rect 39163 34493 39172 34527
rect 39120 34484 39172 34493
rect 39396 34527 39448 34536
rect 39396 34493 39405 34527
rect 39405 34493 39439 34527
rect 39439 34493 39448 34527
rect 39396 34484 39448 34493
rect 37188 34416 37240 34468
rect 22744 34348 22796 34400
rect 27344 34348 27396 34400
rect 28172 34348 28224 34400
rect 33140 34348 33192 34400
rect 37832 34391 37884 34400
rect 37832 34357 37841 34391
rect 37841 34357 37875 34391
rect 37875 34357 37884 34391
rect 37832 34348 37884 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 23388 34144 23440 34196
rect 28080 34144 28132 34196
rect 28356 34144 28408 34196
rect 28540 34187 28592 34196
rect 28540 34153 28549 34187
rect 28549 34153 28583 34187
rect 28583 34153 28592 34187
rect 28540 34144 28592 34153
rect 30472 34187 30524 34196
rect 30472 34153 30481 34187
rect 30481 34153 30515 34187
rect 30515 34153 30524 34187
rect 30472 34144 30524 34153
rect 30840 34144 30892 34196
rect 32312 34144 32364 34196
rect 35716 34144 35768 34196
rect 35992 34187 36044 34196
rect 35992 34153 36001 34187
rect 36001 34153 36035 34187
rect 36035 34153 36044 34187
rect 35992 34144 36044 34153
rect 45744 34144 45796 34196
rect 22468 33983 22520 33992
rect 22468 33949 22477 33983
rect 22477 33949 22511 33983
rect 22511 33949 22520 33983
rect 22468 33940 22520 33949
rect 22744 33983 22796 33992
rect 22744 33949 22778 33983
rect 22778 33949 22796 33983
rect 22744 33940 22796 33949
rect 24952 33940 25004 33992
rect 25320 33983 25372 33992
rect 25320 33949 25329 33983
rect 25329 33949 25363 33983
rect 25363 33949 25372 33983
rect 25320 33940 25372 33949
rect 28264 33940 28316 33992
rect 28908 33940 28960 33992
rect 33784 34076 33836 34128
rect 31576 34008 31628 34060
rect 40408 34051 40460 34060
rect 40408 34017 40417 34051
rect 40417 34017 40451 34051
rect 40451 34017 40460 34051
rect 40408 34008 40460 34017
rect 42800 34076 42852 34128
rect 43260 34008 43312 34060
rect 29644 33940 29696 33992
rect 31392 33940 31444 33992
rect 37280 33940 37332 33992
rect 38108 33983 38160 33992
rect 38108 33949 38142 33983
rect 38142 33949 38160 33983
rect 38108 33940 38160 33949
rect 42064 33940 42116 33992
rect 43076 33940 43128 33992
rect 43168 33940 43220 33992
rect 24400 33804 24452 33856
rect 25136 33847 25188 33856
rect 25136 33813 25145 33847
rect 25145 33813 25179 33847
rect 25179 33813 25188 33847
rect 25136 33804 25188 33813
rect 35348 33872 35400 33924
rect 40040 33872 40092 33924
rect 41328 33872 41380 33924
rect 45376 33983 45428 33992
rect 45376 33949 45385 33983
rect 45385 33949 45419 33983
rect 45419 33949 45428 33983
rect 45376 33940 45428 33949
rect 34060 33804 34112 33856
rect 35808 33847 35860 33856
rect 35808 33813 35833 33847
rect 35833 33813 35860 33847
rect 35808 33804 35860 33813
rect 39028 33804 39080 33856
rect 41236 33804 41288 33856
rect 44456 33872 44508 33924
rect 45192 33872 45244 33924
rect 45652 33940 45704 33992
rect 43720 33847 43772 33856
rect 43720 33813 43729 33847
rect 43729 33813 43763 33847
rect 43763 33813 43772 33847
rect 43720 33804 43772 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 22468 33600 22520 33652
rect 23480 33643 23532 33652
rect 23480 33609 23489 33643
rect 23489 33609 23523 33643
rect 23523 33609 23532 33643
rect 23480 33600 23532 33609
rect 22376 33507 22428 33516
rect 22376 33473 22385 33507
rect 22385 33473 22419 33507
rect 22419 33473 22428 33507
rect 22376 33464 22428 33473
rect 23388 33532 23440 33584
rect 25136 33532 25188 33584
rect 23572 33464 23624 33516
rect 24400 33507 24452 33516
rect 24400 33473 24409 33507
rect 24409 33473 24443 33507
rect 24443 33473 24452 33507
rect 24400 33464 24452 33473
rect 30104 33600 30156 33652
rect 39120 33600 39172 33652
rect 40040 33643 40092 33652
rect 40040 33609 40049 33643
rect 40049 33609 40083 33643
rect 40083 33609 40092 33643
rect 40040 33600 40092 33609
rect 28540 33507 28592 33516
rect 28540 33473 28549 33507
rect 28549 33473 28583 33507
rect 28583 33473 28592 33507
rect 28540 33464 28592 33473
rect 30472 33507 30524 33516
rect 27712 33396 27764 33448
rect 28264 33439 28316 33448
rect 28264 33405 28273 33439
rect 28273 33405 28307 33439
rect 28307 33405 28316 33439
rect 28264 33396 28316 33405
rect 28356 33439 28408 33448
rect 28356 33405 28390 33439
rect 28390 33405 28408 33439
rect 28356 33396 28408 33405
rect 28908 33396 28960 33448
rect 30472 33473 30481 33507
rect 30481 33473 30515 33507
rect 30515 33473 30524 33507
rect 30472 33464 30524 33473
rect 33232 33532 33284 33584
rect 38844 33532 38896 33584
rect 38936 33532 38988 33584
rect 33784 33464 33836 33516
rect 35716 33464 35768 33516
rect 39028 33507 39080 33516
rect 39028 33473 39037 33507
rect 39037 33473 39071 33507
rect 39071 33473 39080 33507
rect 39028 33464 39080 33473
rect 40040 33464 40092 33516
rect 40316 33600 40368 33652
rect 43168 33643 43220 33652
rect 43168 33609 43177 33643
rect 43177 33609 43211 33643
rect 43211 33609 43220 33643
rect 43168 33600 43220 33609
rect 40224 33532 40276 33584
rect 33048 33396 33100 33448
rect 35440 33396 35492 33448
rect 27620 33328 27672 33380
rect 37372 33328 37424 33380
rect 25780 33303 25832 33312
rect 25780 33269 25789 33303
rect 25789 33269 25823 33303
rect 25823 33269 25832 33303
rect 25780 33260 25832 33269
rect 28356 33260 28408 33312
rect 29828 33303 29880 33312
rect 29828 33269 29837 33303
rect 29837 33269 29871 33303
rect 29871 33269 29880 33303
rect 29828 33260 29880 33269
rect 30564 33303 30616 33312
rect 30564 33269 30573 33303
rect 30573 33269 30607 33303
rect 30607 33269 30616 33303
rect 30564 33260 30616 33269
rect 33140 33303 33192 33312
rect 33140 33269 33149 33303
rect 33149 33269 33183 33303
rect 33183 33269 33192 33303
rect 33140 33260 33192 33269
rect 33324 33303 33376 33312
rect 33324 33269 33333 33303
rect 33333 33269 33367 33303
rect 33367 33269 33376 33303
rect 33324 33260 33376 33269
rect 40684 33507 40736 33516
rect 40684 33473 40693 33507
rect 40693 33473 40727 33507
rect 40727 33473 40736 33507
rect 40684 33464 40736 33473
rect 42800 33464 42852 33516
rect 43720 33532 43772 33584
rect 42984 33507 43036 33516
rect 42984 33473 42993 33507
rect 42993 33473 43027 33507
rect 43027 33473 43036 33507
rect 42984 33464 43036 33473
rect 46756 33464 46808 33516
rect 43628 33439 43680 33448
rect 43628 33405 43637 33439
rect 43637 33405 43671 33439
rect 43671 33405 43680 33439
rect 43628 33396 43680 33405
rect 40316 33328 40368 33380
rect 41236 33260 41288 33312
rect 46940 33303 46992 33312
rect 46940 33269 46949 33303
rect 46949 33269 46983 33303
rect 46983 33269 46992 33303
rect 46940 33260 46992 33269
rect 66260 33260 66312 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 24952 33099 25004 33108
rect 24952 33065 24961 33099
rect 24961 33065 24995 33099
rect 24995 33065 25004 33099
rect 24952 33056 25004 33065
rect 27620 33099 27672 33108
rect 27620 33065 27629 33099
rect 27629 33065 27663 33099
rect 27663 33065 27672 33099
rect 27620 33056 27672 33065
rect 28172 33056 28224 33108
rect 33784 33099 33836 33108
rect 33784 33065 33793 33099
rect 33793 33065 33827 33099
rect 33827 33065 33836 33099
rect 33784 33056 33836 33065
rect 35716 33056 35768 33108
rect 42892 33056 42944 33108
rect 43628 33099 43680 33108
rect 43628 33065 43637 33099
rect 43637 33065 43671 33099
rect 43671 33065 43680 33099
rect 43628 33056 43680 33065
rect 23388 32852 23440 32904
rect 26240 32895 26292 32904
rect 26240 32861 26249 32895
rect 26249 32861 26283 32895
rect 26283 32861 26292 32895
rect 26240 32852 26292 32861
rect 25872 32784 25924 32836
rect 29644 32852 29696 32904
rect 29920 32852 29972 32904
rect 31392 32852 31444 32904
rect 32404 32895 32456 32904
rect 32404 32861 32413 32895
rect 32413 32861 32447 32895
rect 32447 32861 32456 32895
rect 32404 32852 32456 32861
rect 35624 32852 35676 32904
rect 37004 32988 37056 33040
rect 67272 32988 67324 33040
rect 37280 32920 37332 32972
rect 46940 32963 46992 32972
rect 37372 32895 37424 32904
rect 26976 32784 27028 32836
rect 27620 32784 27672 32836
rect 22836 32759 22888 32768
rect 22836 32725 22845 32759
rect 22845 32725 22879 32759
rect 22879 32725 22888 32759
rect 22836 32716 22888 32725
rect 27712 32716 27764 32768
rect 28816 32784 28868 32836
rect 32864 32784 32916 32836
rect 33600 32784 33652 32836
rect 37372 32861 37381 32895
rect 37381 32861 37415 32895
rect 37415 32861 37424 32895
rect 37372 32852 37424 32861
rect 37464 32852 37516 32904
rect 46940 32929 46949 32963
rect 46949 32929 46983 32963
rect 46983 32929 46992 32963
rect 46940 32920 46992 32929
rect 66260 32963 66312 32972
rect 66260 32929 66269 32963
rect 66269 32929 66303 32963
rect 66303 32929 66312 32963
rect 66260 32920 66312 32929
rect 42432 32852 42484 32904
rect 42800 32895 42852 32904
rect 42800 32861 42809 32895
rect 42809 32861 42843 32895
rect 42843 32861 42852 32895
rect 42800 32852 42852 32861
rect 43444 32895 43496 32904
rect 43444 32861 43453 32895
rect 43453 32861 43487 32895
rect 43487 32861 43496 32895
rect 43444 32852 43496 32861
rect 44272 32895 44324 32904
rect 44272 32861 44281 32895
rect 44281 32861 44315 32895
rect 44315 32861 44324 32895
rect 44272 32852 44324 32861
rect 46756 32895 46808 32904
rect 46756 32861 46765 32895
rect 46765 32861 46799 32895
rect 46799 32861 46808 32895
rect 46756 32852 46808 32861
rect 36452 32784 36504 32836
rect 65524 32784 65576 32836
rect 66444 32827 66496 32836
rect 66444 32793 66453 32827
rect 66453 32793 66487 32827
rect 66487 32793 66496 32827
rect 66444 32784 66496 32793
rect 68100 32827 68152 32836
rect 68100 32793 68109 32827
rect 68109 32793 68143 32827
rect 68143 32793 68152 32827
rect 68100 32784 68152 32793
rect 28448 32759 28500 32768
rect 28448 32725 28457 32759
rect 28457 32725 28491 32759
rect 28491 32725 28500 32759
rect 28448 32716 28500 32725
rect 29552 32759 29604 32768
rect 29552 32725 29561 32759
rect 29561 32725 29595 32759
rect 29595 32725 29604 32759
rect 29552 32716 29604 32725
rect 30840 32716 30892 32768
rect 34888 32759 34940 32768
rect 34888 32725 34913 32759
rect 34913 32725 34940 32759
rect 34888 32716 34940 32725
rect 36636 32716 36688 32768
rect 38384 32716 38436 32768
rect 39304 32716 39356 32768
rect 43720 32716 43772 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 25320 32512 25372 32564
rect 26240 32512 26292 32564
rect 26976 32555 27028 32564
rect 26976 32521 26985 32555
rect 26985 32521 27019 32555
rect 27019 32521 27028 32555
rect 26976 32512 27028 32521
rect 29644 32512 29696 32564
rect 30104 32555 30156 32564
rect 30104 32521 30113 32555
rect 30113 32521 30147 32555
rect 30147 32521 30156 32555
rect 30104 32512 30156 32521
rect 31392 32555 31444 32564
rect 31392 32521 31401 32555
rect 31401 32521 31435 32555
rect 31435 32521 31444 32555
rect 31392 32512 31444 32521
rect 32404 32555 32456 32564
rect 32404 32521 32413 32555
rect 32413 32521 32447 32555
rect 32447 32521 32456 32555
rect 32404 32512 32456 32521
rect 34888 32512 34940 32564
rect 35808 32512 35860 32564
rect 36452 32555 36504 32564
rect 36452 32521 36461 32555
rect 36461 32521 36495 32555
rect 36495 32521 36504 32555
rect 36452 32512 36504 32521
rect 22836 32444 22888 32496
rect 25780 32444 25832 32496
rect 29552 32444 29604 32496
rect 37372 32444 37424 32496
rect 37648 32444 37700 32496
rect 25504 32419 25556 32428
rect 25504 32385 25513 32419
rect 25513 32385 25547 32419
rect 25547 32385 25556 32419
rect 25504 32376 25556 32385
rect 26056 32376 26108 32428
rect 28448 32376 28500 32428
rect 31300 32376 31352 32428
rect 31852 32376 31904 32428
rect 32312 32419 32364 32428
rect 32312 32385 32321 32419
rect 32321 32385 32355 32419
rect 32355 32385 32364 32419
rect 32312 32376 32364 32385
rect 33784 32376 33836 32428
rect 35440 32376 35492 32428
rect 36636 32419 36688 32428
rect 36636 32385 36645 32419
rect 36645 32385 36679 32419
rect 36679 32385 36688 32419
rect 36636 32376 36688 32385
rect 38384 32419 38436 32428
rect 38384 32385 38393 32419
rect 38393 32385 38427 32419
rect 38427 32385 38436 32419
rect 38384 32376 38436 32385
rect 39396 32444 39448 32496
rect 39488 32444 39540 32496
rect 42616 32444 42668 32496
rect 43720 32444 43772 32496
rect 39304 32419 39356 32428
rect 39304 32385 39313 32419
rect 39313 32385 39347 32419
rect 39347 32385 39356 32419
rect 39304 32376 39356 32385
rect 22376 32351 22428 32360
rect 22376 32317 22385 32351
rect 22385 32317 22419 32351
rect 22419 32317 22428 32351
rect 22376 32308 22428 32317
rect 28724 32351 28776 32360
rect 28724 32317 28733 32351
rect 28733 32317 28767 32351
rect 28767 32317 28776 32351
rect 28724 32308 28776 32317
rect 31944 32308 31996 32360
rect 33600 32351 33652 32360
rect 33600 32317 33609 32351
rect 33609 32317 33643 32351
rect 33643 32317 33652 32351
rect 33600 32308 33652 32317
rect 23020 32172 23072 32224
rect 28264 32240 28316 32292
rect 32956 32240 33008 32292
rect 34428 32351 34480 32360
rect 34428 32317 34462 32351
rect 34462 32317 34480 32351
rect 34428 32308 34480 32317
rect 35348 32308 35400 32360
rect 38292 32351 38344 32360
rect 38292 32317 38301 32351
rect 38301 32317 38335 32351
rect 38335 32317 38344 32351
rect 38292 32308 38344 32317
rect 39580 32419 39632 32428
rect 39580 32385 39614 32419
rect 39614 32385 39632 32419
rect 39580 32376 39632 32385
rect 41144 32376 41196 32428
rect 42432 32376 42484 32428
rect 42708 32419 42760 32428
rect 42708 32385 42717 32419
rect 42717 32385 42751 32419
rect 42751 32385 42760 32419
rect 42708 32376 42760 32385
rect 43076 32376 43128 32428
rect 43628 32376 43680 32428
rect 44364 32419 44416 32428
rect 44364 32385 44373 32419
rect 44373 32385 44407 32419
rect 44407 32385 44416 32419
rect 44364 32376 44416 32385
rect 41328 32308 41380 32360
rect 44548 32419 44600 32428
rect 44548 32385 44557 32419
rect 44557 32385 44591 32419
rect 44591 32385 44600 32419
rect 44548 32376 44600 32385
rect 34060 32283 34112 32292
rect 34060 32249 34069 32283
rect 34069 32249 34103 32283
rect 34103 32249 34112 32283
rect 34060 32240 34112 32249
rect 35900 32215 35952 32224
rect 35900 32181 35909 32215
rect 35909 32181 35943 32215
rect 35943 32181 35952 32215
rect 35900 32172 35952 32181
rect 38108 32215 38160 32224
rect 38108 32181 38117 32215
rect 38117 32181 38151 32215
rect 38151 32181 38160 32215
rect 38108 32172 38160 32181
rect 42064 32240 42116 32292
rect 44640 32308 44692 32360
rect 45560 32444 45612 32496
rect 66444 32512 66496 32564
rect 67272 32376 67324 32428
rect 40684 32215 40736 32224
rect 40684 32181 40693 32215
rect 40693 32181 40727 32215
rect 40727 32181 40736 32215
rect 40684 32172 40736 32181
rect 41328 32172 41380 32224
rect 43352 32172 43404 32224
rect 44364 32172 44416 32224
rect 46756 32172 46808 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 22376 31968 22428 32020
rect 23388 32011 23440 32020
rect 23388 31977 23397 32011
rect 23397 31977 23431 32011
rect 23431 31977 23440 32011
rect 23388 31968 23440 31977
rect 28724 31968 28776 32020
rect 29092 31968 29144 32020
rect 29920 32011 29972 32020
rect 29920 31977 29929 32011
rect 29929 31977 29963 32011
rect 29963 31977 29972 32011
rect 29920 31968 29972 31977
rect 32864 32011 32916 32020
rect 32864 31977 32873 32011
rect 32873 31977 32907 32011
rect 32907 31977 32916 32011
rect 32864 31968 32916 31977
rect 35624 32011 35676 32020
rect 35624 31977 35633 32011
rect 35633 31977 35667 32011
rect 35667 31977 35676 32011
rect 35624 31968 35676 31977
rect 38292 31968 38344 32020
rect 44548 31968 44600 32020
rect 31944 31943 31996 31952
rect 31944 31909 31953 31943
rect 31953 31909 31987 31943
rect 31987 31909 31996 31943
rect 31944 31900 31996 31909
rect 34428 31900 34480 31952
rect 23020 31875 23072 31884
rect 23020 31841 23029 31875
rect 23029 31841 23063 31875
rect 23063 31841 23072 31875
rect 23020 31832 23072 31841
rect 1676 31764 1728 31816
rect 22468 31807 22520 31816
rect 22468 31773 22477 31807
rect 22477 31773 22511 31807
rect 22511 31773 22520 31807
rect 22468 31764 22520 31773
rect 23572 31832 23624 31884
rect 27804 31832 27856 31884
rect 28908 31832 28960 31884
rect 29736 31832 29788 31884
rect 30564 31875 30616 31884
rect 30564 31841 30573 31875
rect 30573 31841 30607 31875
rect 30607 31841 30616 31875
rect 30564 31832 30616 31841
rect 33968 31832 34020 31884
rect 26056 31764 26108 31816
rect 26700 31807 26752 31816
rect 26700 31773 26709 31807
rect 26709 31773 26743 31807
rect 26743 31773 26752 31807
rect 26700 31764 26752 31773
rect 28540 31764 28592 31816
rect 30840 31807 30892 31816
rect 30840 31773 30874 31807
rect 30874 31773 30892 31807
rect 30840 31764 30892 31773
rect 33324 31764 33376 31816
rect 35716 31764 35768 31816
rect 37372 31764 37424 31816
rect 38844 31807 38896 31816
rect 38844 31773 38853 31807
rect 38853 31773 38887 31807
rect 38887 31773 38896 31807
rect 38844 31764 38896 31773
rect 40684 31832 40736 31884
rect 40040 31807 40092 31816
rect 40040 31773 40049 31807
rect 40049 31773 40083 31807
rect 40083 31773 40092 31807
rect 40040 31764 40092 31773
rect 42616 31900 42668 31952
rect 43260 31900 43312 31952
rect 41328 31875 41380 31884
rect 41328 31841 41337 31875
rect 41337 31841 41371 31875
rect 41371 31841 41380 31875
rect 41328 31832 41380 31841
rect 43628 31875 43680 31884
rect 43628 31841 43637 31875
rect 43637 31841 43671 31875
rect 43671 31841 43680 31875
rect 43628 31832 43680 31841
rect 43352 31807 43404 31816
rect 43352 31773 43361 31807
rect 43361 31773 43395 31807
rect 43395 31773 43404 31807
rect 43352 31764 43404 31773
rect 66260 31764 66312 31816
rect 29644 31696 29696 31748
rect 29736 31739 29788 31748
rect 29736 31705 29761 31739
rect 29761 31705 29788 31739
rect 29736 31696 29788 31705
rect 37832 31696 37884 31748
rect 41144 31696 41196 31748
rect 41696 31696 41748 31748
rect 25044 31628 25096 31680
rect 26516 31671 26568 31680
rect 26516 31637 26525 31671
rect 26525 31637 26559 31671
rect 26559 31637 26568 31671
rect 26516 31628 26568 31637
rect 34704 31628 34756 31680
rect 35624 31628 35676 31680
rect 40224 31671 40276 31680
rect 40224 31637 40233 31671
rect 40233 31637 40267 31671
rect 40267 31637 40276 31671
rect 40224 31628 40276 31637
rect 43444 31628 43496 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 22468 31424 22520 31476
rect 23204 31467 23256 31476
rect 23204 31433 23213 31467
rect 23213 31433 23247 31467
rect 23247 31433 23256 31467
rect 23204 31424 23256 31433
rect 26700 31424 26752 31476
rect 27712 31424 27764 31476
rect 39580 31424 39632 31476
rect 41696 31467 41748 31476
rect 41696 31433 41705 31467
rect 41705 31433 41739 31467
rect 41739 31433 41748 31467
rect 41696 31424 41748 31433
rect 26516 31356 26568 31408
rect 1676 31331 1728 31340
rect 1676 31297 1685 31331
rect 1685 31297 1719 31331
rect 1719 31297 1728 31331
rect 1676 31288 1728 31297
rect 25044 31331 25096 31340
rect 2044 31220 2096 31272
rect 2780 31263 2832 31272
rect 2780 31229 2789 31263
rect 2789 31229 2823 31263
rect 2823 31229 2832 31263
rect 2780 31220 2832 31229
rect 25044 31297 25053 31331
rect 25053 31297 25087 31331
rect 25087 31297 25096 31331
rect 25044 31288 25096 31297
rect 27804 31399 27856 31408
rect 27804 31365 27813 31399
rect 27813 31365 27847 31399
rect 27847 31365 27856 31399
rect 27804 31356 27856 31365
rect 34520 31356 34572 31408
rect 35440 31356 35492 31408
rect 35808 31356 35860 31408
rect 38844 31399 38896 31408
rect 38844 31365 38853 31399
rect 38853 31365 38887 31399
rect 38887 31365 38896 31399
rect 38844 31356 38896 31365
rect 39212 31356 39264 31408
rect 32220 31288 32272 31340
rect 32312 31288 32364 31340
rect 34704 31288 34756 31340
rect 35716 31288 35768 31340
rect 37832 31288 37884 31340
rect 38936 31288 38988 31340
rect 40224 31288 40276 31340
rect 42524 31331 42576 31340
rect 42524 31297 42533 31331
rect 42533 31297 42567 31331
rect 42567 31297 42576 31331
rect 42524 31288 42576 31297
rect 42984 31288 43036 31340
rect 43444 31288 43496 31340
rect 44180 31288 44232 31340
rect 66260 31356 66312 31408
rect 43996 31220 44048 31272
rect 65984 31263 66036 31272
rect 65984 31229 65993 31263
rect 65993 31229 66027 31263
rect 66027 31229 66036 31263
rect 65984 31220 66036 31229
rect 67548 31263 67600 31272
rect 67548 31229 67557 31263
rect 67557 31229 67591 31263
rect 67591 31229 67600 31263
rect 67548 31220 67600 31229
rect 26332 31084 26384 31136
rect 26516 31084 26568 31136
rect 28080 31084 28132 31136
rect 28540 31084 28592 31136
rect 31392 31127 31444 31136
rect 31392 31093 31401 31127
rect 31401 31093 31435 31127
rect 31435 31093 31444 31127
rect 31392 31084 31444 31093
rect 33324 31084 33376 31136
rect 35992 31152 36044 31204
rect 35716 31127 35768 31136
rect 35716 31093 35725 31127
rect 35725 31093 35759 31127
rect 35759 31093 35768 31127
rect 35716 31084 35768 31093
rect 36176 31127 36228 31136
rect 36176 31093 36185 31127
rect 36185 31093 36219 31127
rect 36219 31093 36228 31127
rect 36176 31084 36228 31093
rect 37556 31127 37608 31136
rect 37556 31093 37565 31127
rect 37565 31093 37599 31127
rect 37599 31093 37608 31127
rect 37556 31084 37608 31093
rect 39120 31084 39172 31136
rect 43904 31127 43956 31136
rect 43904 31093 43913 31127
rect 43913 31093 43947 31127
rect 43947 31093 43956 31127
rect 43904 31084 43956 31093
rect 44456 31127 44508 31136
rect 44456 31093 44465 31127
rect 44465 31093 44499 31127
rect 44499 31093 44508 31127
rect 44456 31084 44508 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 2044 30923 2096 30932
rect 2044 30889 2053 30923
rect 2053 30889 2087 30923
rect 2087 30889 2096 30923
rect 2044 30880 2096 30889
rect 26332 30880 26384 30932
rect 26792 30880 26844 30932
rect 30472 30880 30524 30932
rect 33140 30880 33192 30932
rect 33416 30923 33468 30932
rect 33416 30889 33425 30923
rect 33425 30889 33459 30923
rect 33459 30889 33468 30923
rect 33416 30880 33468 30889
rect 34704 30923 34756 30932
rect 34704 30889 34713 30923
rect 34713 30889 34747 30923
rect 34747 30889 34756 30923
rect 34704 30880 34756 30889
rect 44180 30923 44232 30932
rect 44180 30889 44189 30923
rect 44189 30889 44223 30923
rect 44223 30889 44232 30923
rect 44180 30880 44232 30889
rect 65984 30880 66036 30932
rect 33232 30744 33284 30796
rect 1952 30719 2004 30728
rect 1952 30685 1961 30719
rect 1961 30685 1995 30719
rect 1995 30685 2004 30719
rect 1952 30676 2004 30685
rect 3332 30676 3384 30728
rect 22468 30719 22520 30728
rect 22468 30685 22477 30719
rect 22477 30685 22511 30719
rect 22511 30685 22520 30719
rect 22468 30676 22520 30685
rect 23204 30719 23256 30728
rect 23204 30685 23213 30719
rect 23213 30685 23247 30719
rect 23247 30685 23256 30719
rect 23204 30676 23256 30685
rect 24584 30719 24636 30728
rect 24584 30685 24593 30719
rect 24593 30685 24627 30719
rect 24627 30685 24636 30719
rect 24584 30676 24636 30685
rect 28540 30719 28592 30728
rect 28540 30685 28549 30719
rect 28549 30685 28583 30719
rect 28583 30685 28592 30719
rect 28540 30676 28592 30685
rect 31116 30719 31168 30728
rect 23480 30608 23532 30660
rect 31116 30685 31125 30719
rect 31125 30685 31159 30719
rect 31159 30685 31168 30719
rect 31116 30676 31168 30685
rect 31392 30719 31444 30728
rect 31392 30685 31426 30719
rect 31426 30685 31444 30719
rect 31392 30676 31444 30685
rect 37556 30787 37608 30796
rect 37556 30753 37565 30787
rect 37565 30753 37599 30787
rect 37599 30753 37608 30787
rect 37556 30744 37608 30753
rect 31760 30608 31812 30660
rect 32312 30608 32364 30660
rect 33324 30608 33376 30660
rect 36176 30676 36228 30728
rect 40040 30676 40092 30728
rect 35348 30608 35400 30660
rect 38200 30608 38252 30660
rect 40132 30608 40184 30660
rect 41144 30676 41196 30728
rect 42708 30676 42760 30728
rect 43996 30719 44048 30728
rect 43996 30685 44005 30719
rect 44005 30685 44039 30719
rect 44039 30685 44048 30719
rect 43996 30676 44048 30685
rect 66812 30676 66864 30728
rect 67548 30719 67600 30728
rect 67548 30685 67557 30719
rect 67557 30685 67591 30719
rect 67591 30685 67600 30719
rect 67548 30676 67600 30685
rect 45468 30608 45520 30660
rect 22100 30540 22152 30592
rect 24400 30583 24452 30592
rect 24400 30549 24409 30583
rect 24409 30549 24443 30583
rect 24443 30549 24452 30583
rect 24400 30540 24452 30549
rect 28356 30583 28408 30592
rect 28356 30549 28365 30583
rect 28365 30549 28399 30583
rect 28399 30549 28408 30583
rect 28356 30540 28408 30549
rect 29644 30583 29696 30592
rect 29644 30549 29653 30583
rect 29653 30549 29687 30583
rect 29687 30549 29696 30583
rect 29644 30540 29696 30549
rect 32496 30583 32548 30592
rect 32496 30549 32505 30583
rect 32505 30549 32539 30583
rect 32539 30549 32548 30583
rect 32496 30540 32548 30549
rect 34520 30540 34572 30592
rect 38844 30540 38896 30592
rect 40776 30583 40828 30592
rect 40776 30549 40785 30583
rect 40785 30549 40819 30583
rect 40819 30549 40828 30583
rect 40776 30540 40828 30549
rect 41420 30583 41472 30592
rect 41420 30549 41429 30583
rect 41429 30549 41463 30583
rect 41463 30549 41472 30583
rect 41420 30540 41472 30549
rect 42984 30540 43036 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 22468 30336 22520 30388
rect 31116 30379 31168 30388
rect 31116 30345 31125 30379
rect 31125 30345 31159 30379
rect 31159 30345 31168 30379
rect 31116 30336 31168 30345
rect 32220 30336 32272 30388
rect 23204 30268 23256 30320
rect 23572 30268 23624 30320
rect 24400 30268 24452 30320
rect 28356 30268 28408 30320
rect 32128 30268 32180 30320
rect 32496 30268 32548 30320
rect 33232 30268 33284 30320
rect 23480 30243 23532 30252
rect 23480 30209 23489 30243
rect 23489 30209 23523 30243
rect 23523 30209 23532 30243
rect 23480 30200 23532 30209
rect 29644 30200 29696 30252
rect 31760 30200 31812 30252
rect 33324 30200 33376 30252
rect 34520 30336 34572 30388
rect 38200 30379 38252 30388
rect 38200 30345 38209 30379
rect 38209 30345 38243 30379
rect 38243 30345 38252 30379
rect 38200 30336 38252 30345
rect 40040 30336 40092 30388
rect 45468 30379 45520 30388
rect 45468 30345 45477 30379
rect 45477 30345 45511 30379
rect 45511 30345 45520 30379
rect 45468 30336 45520 30345
rect 37372 30268 37424 30320
rect 38384 30243 38436 30252
rect 1860 30175 1912 30184
rect 1860 30141 1869 30175
rect 1869 30141 1903 30175
rect 1903 30141 1912 30175
rect 1860 30132 1912 30141
rect 2780 30132 2832 30184
rect 2872 30175 2924 30184
rect 2872 30141 2881 30175
rect 2881 30141 2915 30175
rect 2915 30141 2924 30175
rect 2872 30132 2924 30141
rect 23204 30132 23256 30184
rect 34060 30132 34112 30184
rect 34520 30175 34572 30184
rect 34520 30141 34554 30175
rect 34554 30141 34572 30175
rect 34520 30132 34572 30141
rect 34704 30175 34756 30184
rect 34704 30141 34713 30175
rect 34713 30141 34747 30175
rect 34747 30141 34756 30175
rect 34704 30132 34756 30141
rect 34888 30132 34940 30184
rect 38384 30209 38393 30243
rect 38393 30209 38427 30243
rect 38427 30209 38436 30243
rect 38384 30200 38436 30209
rect 39120 30243 39172 30252
rect 39120 30209 39129 30243
rect 39129 30209 39163 30243
rect 39163 30209 39172 30243
rect 39120 30200 39172 30209
rect 39488 30200 39540 30252
rect 41420 30268 41472 30320
rect 40592 30200 40644 30252
rect 42984 30243 43036 30252
rect 42984 30209 42993 30243
rect 42993 30209 43027 30243
rect 43027 30209 43036 30243
rect 42984 30200 43036 30209
rect 43260 30268 43312 30320
rect 44456 30268 44508 30320
rect 49608 30268 49660 30320
rect 66168 30268 66220 30320
rect 43904 30200 43956 30252
rect 24492 30064 24544 30116
rect 28080 30064 28132 30116
rect 29828 30064 29880 30116
rect 32680 30064 32732 30116
rect 21824 29996 21876 30048
rect 24400 29996 24452 30048
rect 27344 29996 27396 30048
rect 27804 29996 27856 30048
rect 33416 30064 33468 30116
rect 34152 30107 34204 30116
rect 34152 30073 34161 30107
rect 34161 30073 34195 30107
rect 34195 30073 34204 30107
rect 34152 30064 34204 30073
rect 34428 29996 34480 30048
rect 40316 30132 40368 30184
rect 43628 30132 43680 30184
rect 38936 30039 38988 30048
rect 38936 30005 38945 30039
rect 38945 30005 38979 30039
rect 38979 30005 38988 30039
rect 38936 29996 38988 30005
rect 43260 29996 43312 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 1860 29792 1912 29844
rect 2780 29835 2832 29844
rect 2780 29801 2789 29835
rect 2789 29801 2823 29835
rect 2823 29801 2832 29835
rect 2780 29792 2832 29801
rect 23204 29835 23256 29844
rect 23204 29801 23213 29835
rect 23213 29801 23247 29835
rect 23247 29801 23256 29835
rect 23204 29792 23256 29801
rect 24492 29792 24544 29844
rect 24584 29792 24636 29844
rect 27712 29792 27764 29844
rect 34428 29792 34480 29844
rect 35348 29835 35400 29844
rect 35348 29801 35357 29835
rect 35357 29801 35391 29835
rect 35391 29801 35400 29835
rect 35348 29792 35400 29801
rect 38384 29792 38436 29844
rect 21824 29699 21876 29708
rect 21824 29665 21833 29699
rect 21833 29665 21867 29699
rect 21867 29665 21876 29699
rect 21824 29656 21876 29665
rect 24400 29699 24452 29708
rect 24400 29665 24409 29699
rect 24409 29665 24443 29699
rect 24443 29665 24452 29699
rect 24400 29656 24452 29665
rect 4804 29588 4856 29640
rect 22100 29631 22152 29640
rect 22100 29597 22134 29631
rect 22134 29597 22152 29631
rect 22100 29588 22152 29597
rect 23572 29588 23624 29640
rect 25688 29588 25740 29640
rect 25228 29495 25280 29504
rect 25228 29461 25237 29495
rect 25237 29461 25271 29495
rect 25271 29461 25280 29495
rect 25228 29452 25280 29461
rect 26056 29452 26108 29504
rect 26516 29656 26568 29708
rect 32680 29724 32732 29776
rect 34704 29724 34756 29776
rect 34520 29656 34572 29708
rect 43168 29656 43220 29708
rect 27344 29631 27396 29640
rect 27344 29597 27353 29631
rect 27353 29597 27387 29631
rect 27387 29597 27396 29631
rect 27344 29588 27396 29597
rect 29644 29588 29696 29640
rect 29828 29588 29880 29640
rect 31852 29588 31904 29640
rect 35716 29588 35768 29640
rect 37372 29588 37424 29640
rect 38844 29631 38896 29640
rect 38844 29597 38853 29631
rect 38853 29597 38887 29631
rect 38887 29597 38896 29631
rect 38844 29588 38896 29597
rect 30288 29520 30340 29572
rect 27620 29452 27672 29504
rect 29000 29452 29052 29504
rect 39212 29588 39264 29640
rect 40040 29631 40092 29640
rect 40040 29597 40049 29631
rect 40049 29597 40083 29631
rect 40083 29597 40092 29631
rect 40040 29588 40092 29597
rect 40132 29520 40184 29572
rect 40316 29520 40368 29572
rect 43628 29588 43680 29640
rect 46848 29588 46900 29640
rect 31944 29495 31996 29504
rect 31944 29461 31953 29495
rect 31953 29461 31987 29495
rect 31987 29461 31996 29495
rect 31944 29452 31996 29461
rect 38936 29452 38988 29504
rect 39488 29452 39540 29504
rect 40684 29495 40736 29504
rect 40684 29461 40693 29495
rect 40693 29461 40727 29495
rect 40727 29461 40736 29495
rect 40684 29452 40736 29461
rect 44272 29452 44324 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 25228 29180 25280 29232
rect 27804 29248 27856 29300
rect 27896 29248 27948 29300
rect 29000 29291 29052 29300
rect 29000 29257 29009 29291
rect 29009 29257 29043 29291
rect 29043 29257 29052 29291
rect 29000 29248 29052 29257
rect 29644 29291 29696 29300
rect 29644 29257 29653 29291
rect 29653 29257 29687 29291
rect 29687 29257 29696 29291
rect 29644 29248 29696 29257
rect 30288 29291 30340 29300
rect 30288 29257 30297 29291
rect 30297 29257 30331 29291
rect 30331 29257 30340 29291
rect 30288 29248 30340 29257
rect 33968 29291 34020 29300
rect 28080 29155 28132 29164
rect 28080 29121 28089 29155
rect 28089 29121 28123 29155
rect 28123 29121 28132 29155
rect 29644 29155 29696 29164
rect 28080 29112 28132 29121
rect 29644 29121 29653 29155
rect 29653 29121 29687 29155
rect 29687 29121 29696 29155
rect 29644 29112 29696 29121
rect 24676 29087 24728 29096
rect 24676 29053 24685 29087
rect 24685 29053 24719 29087
rect 24719 29053 24728 29087
rect 24676 29044 24728 29053
rect 27436 29044 27488 29096
rect 29828 29044 29880 29096
rect 26056 28951 26108 28960
rect 26056 28917 26065 28951
rect 26065 28917 26099 28951
rect 26099 28917 26108 28951
rect 26056 28908 26108 28917
rect 27804 29019 27856 29028
rect 27804 28985 27813 29019
rect 27813 28985 27847 29019
rect 27847 28985 27856 29019
rect 31944 29112 31996 29164
rect 32128 29155 32180 29164
rect 32128 29121 32137 29155
rect 32137 29121 32171 29155
rect 32171 29121 32180 29155
rect 32128 29112 32180 29121
rect 33968 29257 33977 29291
rect 33977 29257 34011 29291
rect 34011 29257 34020 29291
rect 33968 29248 34020 29257
rect 35256 29291 35308 29300
rect 35256 29257 35281 29291
rect 35281 29257 35308 29291
rect 35256 29248 35308 29257
rect 40592 29291 40644 29300
rect 32496 29044 32548 29096
rect 33140 29087 33192 29096
rect 33140 29053 33174 29087
rect 33174 29053 33192 29087
rect 33140 29044 33192 29053
rect 34704 29044 34756 29096
rect 40592 29257 40601 29291
rect 40601 29257 40635 29291
rect 40635 29257 40644 29291
rect 40592 29248 40644 29257
rect 38108 29180 38160 29232
rect 38200 29155 38252 29164
rect 38200 29121 38209 29155
rect 38209 29121 38243 29155
rect 38243 29121 38252 29155
rect 38200 29112 38252 29121
rect 39304 29155 39356 29164
rect 36544 29044 36596 29096
rect 39304 29121 39313 29155
rect 39313 29121 39347 29155
rect 39347 29121 39356 29155
rect 39304 29112 39356 29121
rect 39488 29155 39540 29164
rect 39488 29121 39497 29155
rect 39497 29121 39531 29155
rect 39531 29121 39540 29155
rect 39488 29112 39540 29121
rect 40224 29112 40276 29164
rect 40776 29155 40828 29164
rect 40776 29121 40785 29155
rect 40785 29121 40819 29155
rect 40819 29121 40828 29155
rect 40776 29112 40828 29121
rect 27804 28976 27856 28985
rect 28816 28908 28868 28960
rect 34152 28976 34204 29028
rect 34704 28908 34756 28960
rect 35992 28976 36044 29028
rect 39304 28976 39356 29028
rect 40224 28976 40276 29028
rect 44364 29248 44416 29300
rect 44272 29223 44324 29232
rect 44272 29189 44281 29223
rect 44281 29189 44315 29223
rect 44315 29189 44324 29223
rect 44272 29180 44324 29189
rect 43260 29155 43312 29164
rect 43260 29121 43269 29155
rect 43269 29121 43303 29155
rect 43303 29121 43312 29155
rect 43260 29112 43312 29121
rect 43720 29112 43772 29164
rect 45928 29087 45980 29096
rect 41512 28976 41564 29028
rect 43720 28976 43772 29028
rect 45928 29053 45937 29087
rect 45937 29053 45971 29087
rect 45971 29053 45980 29087
rect 45928 29044 45980 29053
rect 44180 28976 44232 29028
rect 35900 28951 35952 28960
rect 35900 28917 35909 28951
rect 35909 28917 35943 28951
rect 35943 28917 35952 28951
rect 35900 28908 35952 28917
rect 37924 28951 37976 28960
rect 37924 28917 37933 28951
rect 37933 28917 37967 28951
rect 37967 28917 37976 28951
rect 37924 28908 37976 28917
rect 39120 28908 39172 28960
rect 42892 28908 42944 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 24676 28704 24728 28756
rect 25688 28747 25740 28756
rect 25688 28713 25697 28747
rect 25697 28713 25731 28747
rect 25731 28713 25740 28747
rect 25688 28704 25740 28713
rect 29092 28704 29144 28756
rect 34704 28704 34756 28756
rect 36544 28747 36596 28756
rect 36544 28713 36553 28747
rect 36553 28713 36587 28747
rect 36587 28713 36596 28747
rect 36544 28704 36596 28713
rect 44180 28747 44232 28756
rect 44180 28713 44189 28747
rect 44189 28713 44223 28747
rect 44223 28713 44232 28747
rect 44180 28704 44232 28713
rect 26056 28568 26108 28620
rect 31760 28568 31812 28620
rect 33048 28568 33100 28620
rect 40408 28568 40460 28620
rect 25504 28543 25556 28552
rect 25504 28509 25513 28543
rect 25513 28509 25547 28543
rect 25547 28509 25556 28543
rect 25504 28500 25556 28509
rect 24952 28432 25004 28484
rect 29644 28500 29696 28552
rect 31852 28500 31904 28552
rect 35164 28543 35216 28552
rect 35164 28509 35173 28543
rect 35173 28509 35207 28543
rect 35207 28509 35216 28543
rect 35164 28500 35216 28509
rect 35900 28500 35952 28552
rect 42892 28500 42944 28552
rect 37924 28432 37976 28484
rect 40868 28432 40920 28484
rect 26332 28407 26384 28416
rect 26332 28373 26341 28407
rect 26341 28373 26375 28407
rect 26375 28373 26384 28407
rect 26332 28364 26384 28373
rect 30196 28364 30248 28416
rect 31392 28364 31444 28416
rect 31668 28364 31720 28416
rect 38200 28364 38252 28416
rect 41052 28364 41104 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 31668 28160 31720 28212
rect 35164 28160 35216 28212
rect 40868 28203 40920 28212
rect 40868 28169 40877 28203
rect 40877 28169 40911 28203
rect 40911 28169 40920 28203
rect 40868 28160 40920 28169
rect 25504 28092 25556 28144
rect 27620 28092 27672 28144
rect 28816 28135 28868 28144
rect 28816 28101 28825 28135
rect 28825 28101 28859 28135
rect 28859 28101 28868 28135
rect 28816 28092 28868 28101
rect 29736 28092 29788 28144
rect 30196 28067 30248 28076
rect 30196 28033 30205 28067
rect 30205 28033 30239 28067
rect 30239 28033 30248 28067
rect 30196 28024 30248 28033
rect 31208 28024 31260 28076
rect 34796 28024 34848 28076
rect 23204 27999 23256 28008
rect 23204 27965 23213 27999
rect 23213 27965 23247 27999
rect 23247 27965 23256 27999
rect 23204 27956 23256 27965
rect 13820 27888 13872 27940
rect 26516 27956 26568 28008
rect 27436 27956 27488 28008
rect 28908 27956 28960 28008
rect 26608 27820 26660 27872
rect 28356 27863 28408 27872
rect 28356 27829 28365 27863
rect 28365 27829 28399 27863
rect 28399 27829 28408 27863
rect 28356 27820 28408 27829
rect 29092 27888 29144 27940
rect 29184 27863 29236 27872
rect 29184 27829 29193 27863
rect 29193 27829 29227 27863
rect 29227 27829 29236 27863
rect 29184 27820 29236 27829
rect 34336 27999 34388 28008
rect 34336 27965 34345 27999
rect 34345 27965 34379 27999
rect 34379 27965 34388 27999
rect 34336 27956 34388 27965
rect 34520 27956 34572 28008
rect 35624 28024 35676 28076
rect 40408 28092 40460 28144
rect 39120 28067 39172 28076
rect 39120 28033 39154 28067
rect 39154 28033 39172 28067
rect 39120 28024 39172 28033
rect 40040 28024 40092 28076
rect 41052 28024 41104 28076
rect 44364 28092 44416 28144
rect 41512 28067 41564 28076
rect 40684 27956 40736 28008
rect 41512 28033 41521 28067
rect 41521 28033 41555 28067
rect 41555 28033 41564 28067
rect 41512 28024 41564 28033
rect 31760 27888 31812 27940
rect 33232 27863 33284 27872
rect 33232 27829 33241 27863
rect 33241 27829 33275 27863
rect 33275 27829 33284 27863
rect 33232 27820 33284 27829
rect 40224 27863 40276 27872
rect 40224 27829 40233 27863
rect 40233 27829 40267 27863
rect 40267 27829 40276 27863
rect 40224 27820 40276 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 23204 27659 23256 27668
rect 23204 27625 23213 27659
rect 23213 27625 23247 27659
rect 23247 27625 23256 27659
rect 23204 27616 23256 27625
rect 27620 27616 27672 27668
rect 31208 27659 31260 27668
rect 31208 27625 31217 27659
rect 31217 27625 31251 27659
rect 31251 27625 31260 27659
rect 31208 27616 31260 27625
rect 34060 27591 34112 27600
rect 34060 27557 34069 27591
rect 34069 27557 34103 27591
rect 34103 27557 34112 27591
rect 34060 27548 34112 27557
rect 26148 27523 26200 27532
rect 26148 27489 26157 27523
rect 26157 27489 26191 27523
rect 26191 27489 26200 27523
rect 26148 27480 26200 27489
rect 28816 27480 28868 27532
rect 30012 27480 30064 27532
rect 24308 27412 24360 27464
rect 26976 27455 27028 27464
rect 26976 27421 26985 27455
rect 26985 27421 27019 27455
rect 27019 27421 27028 27455
rect 26976 27412 27028 27421
rect 29184 27412 29236 27464
rect 30472 27455 30524 27464
rect 24584 27387 24636 27396
rect 24584 27353 24593 27387
rect 24593 27353 24627 27387
rect 24627 27353 24636 27387
rect 24584 27344 24636 27353
rect 27528 27344 27580 27396
rect 27620 27344 27672 27396
rect 30472 27421 30481 27455
rect 30481 27421 30515 27455
rect 30515 27421 30524 27455
rect 30472 27412 30524 27421
rect 31392 27455 31444 27464
rect 31392 27421 31401 27455
rect 31401 27421 31435 27455
rect 31435 27421 31444 27455
rect 31392 27412 31444 27421
rect 32680 27455 32732 27464
rect 32680 27421 32689 27455
rect 32689 27421 32723 27455
rect 32723 27421 32732 27455
rect 32680 27412 32732 27421
rect 33232 27412 33284 27464
rect 34520 27480 34572 27532
rect 34796 27548 34848 27600
rect 33968 27412 34020 27464
rect 34336 27412 34388 27464
rect 34244 27344 34296 27396
rect 38476 27548 38528 27600
rect 40224 27548 40276 27600
rect 37372 27387 37424 27396
rect 37372 27353 37381 27387
rect 37381 27353 37415 27387
rect 37415 27353 37424 27387
rect 37372 27344 37424 27353
rect 28724 27276 28776 27328
rect 28908 27276 28960 27328
rect 29736 27319 29788 27328
rect 29736 27285 29745 27319
rect 29745 27285 29779 27319
rect 29779 27285 29788 27319
rect 29736 27276 29788 27285
rect 30656 27319 30708 27328
rect 30656 27285 30665 27319
rect 30665 27285 30699 27319
rect 30699 27285 30708 27319
rect 30656 27276 30708 27285
rect 32864 27276 32916 27328
rect 40868 27455 40920 27464
rect 40868 27421 40877 27455
rect 40877 27421 40911 27455
rect 40911 27421 40920 27455
rect 40868 27412 40920 27421
rect 41512 27276 41564 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 24584 27072 24636 27124
rect 26516 27072 26568 27124
rect 26976 27072 27028 27124
rect 28724 27072 28776 27124
rect 30012 27115 30064 27124
rect 26608 27004 26660 27056
rect 24308 26936 24360 26988
rect 26332 26936 26384 26988
rect 27620 26936 27672 26988
rect 29736 27004 29788 27056
rect 30012 27081 30021 27115
rect 30021 27081 30055 27115
rect 30055 27081 30064 27115
rect 30012 27072 30064 27081
rect 32680 27115 32732 27124
rect 32680 27081 32689 27115
rect 32689 27081 32723 27115
rect 32723 27081 32732 27115
rect 32680 27072 32732 27081
rect 34244 27004 34296 27056
rect 28908 26979 28960 26988
rect 28908 26945 28942 26979
rect 28942 26945 28960 26979
rect 28908 26936 28960 26945
rect 30656 26936 30708 26988
rect 33140 26936 33192 26988
rect 33968 26979 34020 26988
rect 33968 26945 33977 26979
rect 33977 26945 34011 26979
rect 34011 26945 34020 26979
rect 33968 26936 34020 26945
rect 35532 27072 35584 27124
rect 37372 27115 37424 27124
rect 37372 27081 37381 27115
rect 37381 27081 37415 27115
rect 37415 27081 37424 27115
rect 37372 27072 37424 27081
rect 34704 26936 34756 26988
rect 35440 26936 35492 26988
rect 40040 26979 40092 26988
rect 24216 26732 24268 26784
rect 35624 26732 35676 26784
rect 40040 26945 40049 26979
rect 40049 26945 40083 26979
rect 40083 26945 40092 26979
rect 40040 26936 40092 26945
rect 40316 26868 40368 26920
rect 38844 26800 38896 26852
rect 45744 26732 45796 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 27528 26571 27580 26580
rect 27528 26537 27537 26571
rect 27537 26537 27571 26571
rect 27571 26537 27580 26571
rect 27528 26528 27580 26537
rect 34704 26571 34756 26580
rect 24308 26460 24360 26512
rect 32956 26435 33008 26444
rect 32956 26401 32965 26435
rect 32965 26401 32999 26435
rect 32999 26401 33008 26435
rect 32956 26392 33008 26401
rect 34704 26537 34713 26571
rect 34713 26537 34747 26571
rect 34747 26537 34756 26571
rect 34704 26528 34756 26537
rect 35440 26571 35492 26580
rect 35440 26537 35449 26571
rect 35449 26537 35483 26571
rect 35483 26537 35492 26571
rect 35440 26528 35492 26537
rect 40316 26571 40368 26580
rect 40316 26537 40325 26571
rect 40325 26537 40359 26571
rect 40359 26537 40368 26571
rect 40316 26528 40368 26537
rect 1676 26324 1728 26376
rect 3056 26324 3108 26376
rect 28356 26324 28408 26376
rect 31116 26367 31168 26376
rect 31116 26333 31125 26367
rect 31125 26333 31159 26367
rect 31159 26333 31168 26367
rect 31116 26324 31168 26333
rect 32864 26324 32916 26376
rect 33140 26367 33192 26376
rect 33140 26333 33149 26367
rect 33149 26333 33183 26367
rect 33183 26333 33192 26367
rect 33140 26324 33192 26333
rect 33784 26324 33836 26376
rect 35624 26367 35676 26376
rect 35624 26333 35633 26367
rect 35633 26333 35667 26367
rect 35667 26333 35676 26367
rect 35624 26324 35676 26333
rect 40868 26392 40920 26444
rect 41236 26392 41288 26444
rect 41512 26435 41564 26444
rect 41512 26401 41521 26435
rect 41521 26401 41555 26435
rect 41555 26401 41564 26435
rect 41512 26392 41564 26401
rect 32128 26256 32180 26308
rect 43168 26299 43220 26308
rect 43168 26265 43177 26299
rect 43177 26265 43211 26299
rect 43211 26265 43220 26299
rect 43168 26256 43220 26265
rect 33324 26231 33376 26240
rect 33324 26197 33333 26231
rect 33333 26197 33367 26231
rect 33367 26197 33376 26231
rect 33324 26188 33376 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 31116 26027 31168 26036
rect 31116 25993 31125 26027
rect 31125 25993 31159 26027
rect 31159 25993 31168 26027
rect 31116 25984 31168 25993
rect 32128 26027 32180 26036
rect 32128 25993 32137 26027
rect 32137 25993 32171 26027
rect 32171 25993 32180 26027
rect 32128 25984 32180 25993
rect 34796 25984 34848 26036
rect 30656 25916 30708 25968
rect 1676 25891 1728 25900
rect 1676 25857 1685 25891
rect 1685 25857 1719 25891
rect 1719 25857 1728 25891
rect 1676 25848 1728 25857
rect 31392 25916 31444 25968
rect 33784 25916 33836 25968
rect 33324 25848 33376 25900
rect 33968 25891 34020 25900
rect 33968 25857 34002 25891
rect 34002 25857 34020 25891
rect 33968 25848 34020 25857
rect 2320 25780 2372 25832
rect 2780 25823 2832 25832
rect 2780 25789 2789 25823
rect 2789 25789 2823 25823
rect 2823 25789 2832 25823
rect 2780 25780 2832 25789
rect 33692 25823 33744 25832
rect 33692 25789 33701 25823
rect 33701 25789 33735 25823
rect 33735 25789 33744 25823
rect 33692 25780 33744 25789
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 2320 25483 2372 25492
rect 2320 25449 2329 25483
rect 2329 25449 2363 25483
rect 2363 25449 2372 25483
rect 2320 25440 2372 25449
rect 33692 25440 33744 25492
rect 32496 25347 32548 25356
rect 32496 25313 32505 25347
rect 32505 25313 32539 25347
rect 32539 25313 32548 25347
rect 32496 25304 32548 25313
rect 3424 25236 3476 25288
rect 33140 25236 33192 25288
rect 33784 25279 33836 25288
rect 33784 25245 33793 25279
rect 33793 25245 33827 25279
rect 33827 25245 33836 25279
rect 33784 25236 33836 25245
rect 34796 25279 34848 25288
rect 34796 25245 34805 25279
rect 34805 25245 34839 25279
rect 34839 25245 34848 25279
rect 34796 25236 34848 25245
rect 32404 25100 32456 25152
rect 35072 25143 35124 25152
rect 35072 25109 35081 25143
rect 35081 25109 35115 25143
rect 35115 25109 35124 25143
rect 35072 25100 35124 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 33968 24896 34020 24948
rect 1860 24803 1912 24812
rect 1860 24769 1869 24803
rect 1869 24769 1903 24803
rect 1903 24769 1912 24803
rect 1860 24760 1912 24769
rect 5264 24760 5316 24812
rect 31392 24803 31444 24812
rect 31392 24769 31401 24803
rect 31401 24769 31435 24803
rect 31435 24769 31444 24803
rect 31392 24760 31444 24769
rect 32220 24760 32272 24812
rect 35072 24760 35124 24812
rect 2044 24556 2096 24608
rect 3424 24599 3476 24608
rect 3424 24565 3433 24599
rect 3433 24565 3467 24599
rect 3467 24565 3476 24599
rect 3424 24556 3476 24565
rect 20720 24556 20772 24608
rect 32496 24556 32548 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 32220 24395 32272 24404
rect 32220 24361 32229 24395
rect 32229 24361 32263 24395
rect 32263 24361 32272 24395
rect 32220 24352 32272 24361
rect 3424 24284 3476 24336
rect 2044 24216 2096 24268
rect 2780 24259 2832 24268
rect 2780 24225 2789 24259
rect 2789 24225 2823 24259
rect 2823 24225 2832 24259
rect 2780 24216 2832 24225
rect 32404 24191 32456 24200
rect 32404 24157 32413 24191
rect 32413 24157 32447 24191
rect 32447 24157 32456 24191
rect 32404 24148 32456 24157
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 66260 23468 66312 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 66260 23171 66312 23180
rect 66260 23137 66269 23171
rect 66269 23137 66303 23171
rect 66303 23137 66312 23171
rect 66260 23128 66312 23137
rect 68100 23171 68152 23180
rect 68100 23137 68109 23171
rect 68109 23137 68143 23171
rect 68143 23137 68152 23171
rect 68100 23128 68152 23137
rect 66444 23035 66496 23044
rect 66444 23001 66453 23035
rect 66453 23001 66487 23035
rect 66487 23001 66496 23035
rect 66444 22992 66496 23001
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 66444 22720 66496 22772
rect 67180 22627 67232 22636
rect 67180 22593 67189 22627
rect 67189 22593 67223 22627
rect 67223 22593 67232 22627
rect 67180 22584 67232 22593
rect 1768 22559 1820 22568
rect 1768 22525 1777 22559
rect 1777 22525 1811 22559
rect 1811 22525 1820 22559
rect 1768 22516 1820 22525
rect 2596 22516 2648 22568
rect 2780 22559 2832 22568
rect 2780 22525 2789 22559
rect 2789 22525 2823 22559
rect 2823 22525 2832 22559
rect 2780 22516 2832 22525
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 1768 22176 1820 22228
rect 2596 22219 2648 22228
rect 2596 22185 2605 22219
rect 2605 22185 2639 22219
rect 2639 22185 2648 22219
rect 2596 22176 2648 22185
rect 66260 22108 66312 22160
rect 4620 21972 4672 22024
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 65984 21607 66036 21616
rect 65984 21573 65993 21607
rect 65993 21573 66027 21607
rect 66027 21573 66036 21607
rect 65984 21564 66036 21573
rect 1860 21539 1912 21548
rect 1860 21505 1869 21539
rect 1869 21505 1903 21539
rect 1903 21505 1912 21539
rect 1860 21496 1912 21505
rect 66260 21428 66312 21480
rect 67548 21471 67600 21480
rect 67548 21437 67557 21471
rect 67557 21437 67591 21471
rect 67591 21437 67600 21471
rect 67548 21428 67600 21437
rect 19156 21292 19208 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 67824 18751 67876 18760
rect 67824 18717 67833 18751
rect 67833 18717 67867 18751
rect 67867 18717 67876 18751
rect 67824 18708 67876 18717
rect 68008 18615 68060 18624
rect 68008 18581 68017 18615
rect 68017 18581 68051 18615
rect 68051 18581 68060 18615
rect 68008 18572 68060 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 28724 18300 28776 18352
rect 68008 18232 68060 18284
rect 27436 18164 27488 18216
rect 3976 18096 4028 18148
rect 36912 18028 36964 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 65800 17620 65852 17672
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 67732 17212 67784 17264
rect 65800 17187 65852 17196
rect 65800 17153 65809 17187
rect 65809 17153 65843 17187
rect 65843 17153 65852 17187
rect 65800 17144 65852 17153
rect 67548 17119 67600 17128
rect 67548 17085 67557 17119
rect 67557 17085 67591 17119
rect 67591 17085 67600 17119
rect 67548 17076 67600 17085
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 66720 16600 66772 16652
rect 43168 16532 43220 16584
rect 66168 16532 66220 16584
rect 67732 16396 67784 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 2044 16031 2096 16040
rect 2044 15997 2053 16031
rect 2053 15997 2087 16031
rect 2087 15997 2096 16031
rect 2044 15988 2096 15997
rect 2872 15988 2924 16040
rect 2964 16031 3016 16040
rect 2964 15997 2973 16031
rect 2973 15997 3007 16031
rect 3007 15997 3016 16031
rect 2964 15988 3016 15997
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 2044 15648 2096 15700
rect 2872 15691 2924 15700
rect 2872 15657 2881 15691
rect 2881 15657 2915 15691
rect 2915 15657 2924 15691
rect 2872 15648 2924 15657
rect 2872 15444 2924 15496
rect 4712 15444 4764 15496
rect 67272 15444 67324 15496
rect 66260 15308 66312 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 66260 15036 66312 15088
rect 67364 14900 67416 14952
rect 67548 14943 67600 14952
rect 67548 14909 67557 14943
rect 67557 14909 67591 14943
rect 67591 14909 67600 14943
rect 67548 14900 67600 14909
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 67364 14560 67416 14612
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 1584 13268 1636 13320
rect 67824 13311 67876 13320
rect 67824 13277 67833 13311
rect 67833 13277 67867 13311
rect 67867 13277 67876 13311
rect 67824 13268 67876 13277
rect 68008 13175 68060 13184
rect 68008 13141 68017 13175
rect 68017 13141 68051 13175
rect 68051 13141 68060 13175
rect 68008 13132 68060 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 1584 12835 1636 12844
rect 1584 12801 1593 12835
rect 1593 12801 1627 12835
rect 1627 12801 1636 12835
rect 1584 12792 1636 12801
rect 32128 12835 32180 12844
rect 32128 12801 32137 12835
rect 32137 12801 32171 12835
rect 32171 12801 32180 12835
rect 32128 12792 32180 12801
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 2780 12724 2832 12733
rect 31944 12724 31996 12776
rect 68008 12724 68060 12776
rect 22560 12588 22612 12640
rect 32404 12631 32456 12640
rect 32404 12597 32413 12631
rect 32413 12597 32447 12631
rect 32447 12597 32456 12631
rect 32404 12588 32456 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 1768 12384 1820 12436
rect 2412 12180 2464 12232
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 67640 7871 67692 7880
rect 67640 7837 67649 7871
rect 67649 7837 67683 7871
rect 67683 7837 67692 7871
rect 67640 7828 67692 7837
rect 1860 7803 1912 7812
rect 1860 7769 1869 7803
rect 1869 7769 1903 7803
rect 1903 7769 1912 7803
rect 1860 7760 1912 7769
rect 19984 7760 20036 7812
rect 17592 7692 17644 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 65800 6740 65852 6792
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 65800 6307 65852 6316
rect 65800 6273 65809 6307
rect 65809 6273 65843 6307
rect 65843 6273 65852 6307
rect 65800 6264 65852 6273
rect 65984 6239 66036 6248
rect 65984 6205 65993 6239
rect 65993 6205 66027 6239
rect 66027 6205 66036 6239
rect 65984 6196 66036 6205
rect 67548 6239 67600 6248
rect 67548 6205 67557 6239
rect 67557 6205 67591 6239
rect 67591 6205 67600 6239
rect 67548 6196 67600 6205
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 65984 5856 66036 5908
rect 2780 5652 2832 5704
rect 66444 5695 66496 5704
rect 66444 5661 66453 5695
rect 66453 5661 66487 5695
rect 66487 5661 66496 5695
rect 66444 5652 66496 5661
rect 67272 5652 67324 5704
rect 66996 5559 67048 5568
rect 66996 5525 67005 5559
rect 67005 5525 67039 5559
rect 67039 5525 67048 5559
rect 66996 5516 67048 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 66996 5244 67048 5296
rect 66444 5108 66496 5160
rect 67548 5151 67600 5160
rect 67548 5117 67557 5151
rect 67557 5117 67591 5151
rect 67591 5117 67600 5151
rect 67548 5108 67600 5117
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 24124 4564 24176 4616
rect 66904 4607 66956 4616
rect 66904 4573 66913 4607
rect 66913 4573 66947 4607
rect 66947 4573 66956 4607
rect 66904 4564 66956 4573
rect 67272 4564 67324 4616
rect 6368 4496 6420 4548
rect 10232 4496 10284 4548
rect 67456 4471 67508 4480
rect 67456 4437 67465 4471
rect 67465 4437 67499 4471
rect 67499 4437 67508 4471
rect 67456 4428 67508 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 6368 4088 6420 4140
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 34612 4088 34664 4140
rect 36084 4088 36136 4140
rect 45744 4131 45796 4140
rect 45744 4097 45753 4131
rect 45753 4097 45787 4131
rect 45787 4097 45796 4131
rect 45744 4088 45796 4097
rect 41236 4020 41288 4072
rect 45928 4020 45980 4072
rect 1584 3884 1636 3936
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 4620 3884 4672 3893
rect 5172 3927 5224 3936
rect 5172 3893 5181 3927
rect 5181 3893 5215 3927
rect 5215 3893 5224 3927
rect 5172 3884 5224 3893
rect 6828 3884 6880 3936
rect 46388 3884 46440 3936
rect 60648 3884 60700 3936
rect 62120 3884 62172 3936
rect 67456 4020 67508 4072
rect 68928 4020 68980 4072
rect 66904 3952 66956 4004
rect 67180 3884 67232 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 664 3680 716 3732
rect 3148 3612 3200 3664
rect 4620 3544 4672 3596
rect 47676 3612 47728 3664
rect 10968 3587 11020 3596
rect 1952 3519 2004 3528
rect 1952 3485 1961 3519
rect 1961 3485 1995 3519
rect 1995 3485 2004 3519
rect 1952 3476 2004 3485
rect 3884 3476 3936 3528
rect 5172 3408 5224 3460
rect 6644 3408 6696 3460
rect 1768 3340 1820 3392
rect 6552 3340 6604 3392
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 10416 3519 10468 3528
rect 10416 3485 10425 3519
rect 10425 3485 10459 3519
rect 10459 3485 10468 3519
rect 10416 3476 10468 3485
rect 10600 3451 10652 3460
rect 10600 3417 10609 3451
rect 10609 3417 10643 3451
rect 10643 3417 10652 3451
rect 10600 3408 10652 3417
rect 19340 3476 19392 3528
rect 23112 3544 23164 3596
rect 46388 3587 46440 3596
rect 23848 3476 23900 3528
rect 38108 3476 38160 3528
rect 46388 3553 46397 3587
rect 46397 3553 46431 3587
rect 46431 3553 46440 3587
rect 46388 3544 46440 3553
rect 47032 3587 47084 3596
rect 47032 3553 47041 3587
rect 47041 3553 47075 3587
rect 47075 3553 47084 3587
rect 47032 3544 47084 3553
rect 62120 3587 62172 3596
rect 62120 3553 62129 3587
rect 62129 3553 62163 3587
rect 62163 3553 62172 3587
rect 62120 3544 62172 3553
rect 62488 3587 62540 3596
rect 62488 3553 62497 3587
rect 62497 3553 62531 3587
rect 62531 3553 62540 3587
rect 62488 3544 62540 3553
rect 46204 3519 46256 3528
rect 46204 3485 46213 3519
rect 46213 3485 46247 3519
rect 46247 3485 46256 3519
rect 46204 3476 46256 3485
rect 50896 3476 50948 3528
rect 51724 3476 51776 3528
rect 59728 3476 59780 3528
rect 25596 3408 25648 3460
rect 43812 3408 43864 3460
rect 65800 3476 65852 3528
rect 67364 3476 67416 3528
rect 62120 3408 62172 3460
rect 22100 3383 22152 3392
rect 22100 3349 22109 3383
rect 22109 3349 22143 3383
rect 22143 3349 22152 3383
rect 22100 3340 22152 3349
rect 24492 3340 24544 3392
rect 26148 3340 26200 3392
rect 44824 3340 44876 3392
rect 60832 3383 60884 3392
rect 60832 3349 60841 3383
rect 60841 3349 60875 3383
rect 60875 3349 60884 3383
rect 60832 3340 60884 3349
rect 65984 3340 66036 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 1952 3136 2004 3188
rect 37280 3136 37332 3188
rect 1768 3111 1820 3120
rect 1768 3077 1777 3111
rect 1777 3077 1811 3111
rect 1811 3077 1820 3111
rect 1768 3068 1820 3077
rect 6828 3111 6880 3120
rect 6828 3077 6837 3111
rect 6837 3077 6871 3111
rect 6871 3077 6880 3111
rect 6828 3068 6880 3077
rect 10600 3111 10652 3120
rect 10600 3077 10609 3111
rect 10609 3077 10643 3111
rect 10643 3077 10652 3111
rect 10600 3068 10652 3077
rect 22100 3111 22152 3120
rect 22100 3077 22109 3111
rect 22109 3077 22143 3111
rect 22143 3077 22152 3111
rect 22100 3068 22152 3077
rect 44824 3111 44876 3120
rect 44824 3077 44833 3111
rect 44833 3077 44867 3111
rect 44867 3077 44876 3111
rect 44824 3068 44876 3077
rect 60832 3111 60884 3120
rect 60832 3077 60841 3111
rect 60841 3077 60875 3111
rect 60875 3077 60884 3111
rect 60832 3068 60884 3077
rect 65984 3111 66036 3120
rect 65984 3077 65993 3111
rect 65993 3077 66027 3111
rect 66027 3077 66036 3111
rect 65984 3068 66036 3077
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 10232 3043 10284 3052
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 19340 3043 19392 3052
rect 2780 2975 2832 2984
rect 2780 2941 2789 2975
rect 2789 2941 2823 2975
rect 2823 2941 2832 2975
rect 2780 2932 2832 2941
rect 3516 2932 3568 2984
rect 7104 2975 7156 2984
rect 2872 2864 2924 2916
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 19340 3009 19349 3043
rect 19349 3009 19383 3043
rect 19383 3009 19392 3043
rect 19340 3000 19392 3009
rect 33416 3043 33468 3052
rect 33416 3009 33425 3043
rect 33425 3009 33459 3043
rect 33459 3009 33468 3043
rect 33416 3000 33468 3009
rect 38108 3043 38160 3052
rect 38108 3009 38117 3043
rect 38117 3009 38151 3043
rect 38151 3009 38160 3043
rect 38108 3000 38160 3009
rect 60648 3043 60700 3052
rect 60648 3009 60657 3043
rect 60657 3009 60691 3043
rect 60691 3009 60700 3043
rect 60648 3000 60700 3009
rect 65800 3043 65852 3052
rect 65800 3009 65809 3043
rect 65809 3009 65843 3043
rect 65843 3009 65852 3043
rect 65800 3000 65852 3009
rect 19524 2975 19576 2984
rect 19524 2941 19533 2975
rect 19533 2941 19567 2975
rect 19567 2941 19576 2975
rect 19524 2932 19576 2941
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 22744 2932 22796 2984
rect 22560 2864 22612 2916
rect 34612 2932 34664 2984
rect 34796 2975 34848 2984
rect 34796 2941 34805 2975
rect 34805 2941 34839 2975
rect 34839 2941 34848 2975
rect 34796 2932 34848 2941
rect 38292 2975 38344 2984
rect 38292 2941 38301 2975
rect 38301 2941 38335 2975
rect 38335 2941 38344 2975
rect 38292 2932 38344 2941
rect 38660 2975 38712 2984
rect 38660 2941 38669 2975
rect 38669 2941 38703 2975
rect 38703 2941 38712 2975
rect 38660 2932 38712 2941
rect 45100 2975 45152 2984
rect 45100 2941 45109 2975
rect 45109 2941 45143 2975
rect 45143 2941 45152 2975
rect 45100 2932 45152 2941
rect 61200 2975 61252 2984
rect 61200 2941 61209 2975
rect 61209 2941 61243 2975
rect 61243 2941 61252 2975
rect 61200 2932 61252 2941
rect 69572 2932 69624 2984
rect 67088 2864 67140 2916
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 3516 2592 3568 2644
rect 3976 2635 4028 2644
rect 3976 2601 3985 2635
rect 3985 2601 4019 2635
rect 4019 2601 4028 2635
rect 3976 2592 4028 2601
rect 10416 2592 10468 2644
rect 17684 2635 17736 2644
rect 17684 2601 17693 2635
rect 17693 2601 17727 2635
rect 17727 2601 17736 2635
rect 17684 2592 17736 2601
rect 19524 2635 19576 2644
rect 19524 2601 19533 2635
rect 19533 2601 19567 2635
rect 19567 2601 19576 2635
rect 19524 2592 19576 2601
rect 22744 2635 22796 2644
rect 22744 2601 22753 2635
rect 22753 2601 22787 2635
rect 22787 2601 22796 2635
rect 22744 2592 22796 2601
rect 32312 2635 32364 2644
rect 32312 2601 32321 2635
rect 32321 2601 32355 2635
rect 32355 2601 32364 2635
rect 32312 2592 32364 2601
rect 34612 2592 34664 2644
rect 38292 2592 38344 2644
rect 46204 2592 46256 2644
rect 62120 2635 62172 2644
rect 62120 2601 62129 2635
rect 62129 2601 62163 2635
rect 62163 2601 62172 2635
rect 62120 2592 62172 2601
rect 5816 2524 5868 2576
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 25412 2524 25464 2576
rect 25964 2524 26016 2576
rect 2412 2431 2464 2440
rect 2412 2397 2421 2431
rect 2421 2397 2455 2431
rect 2455 2397 2464 2431
rect 2412 2388 2464 2397
rect 3240 2388 3292 2440
rect 17408 2388 17460 2440
rect 25320 2456 25372 2508
rect 27436 2499 27488 2508
rect 21272 2388 21324 2440
rect 27068 2388 27120 2440
rect 27436 2465 27445 2499
rect 27445 2465 27479 2499
rect 27479 2465 27488 2499
rect 27436 2456 27488 2465
rect 33416 2456 33468 2508
rect 28356 2388 28408 2440
rect 32220 2388 32272 2440
rect 37280 2388 37332 2440
rect 20904 2320 20956 2372
rect 20812 2252 20864 2304
rect 32128 2252 32180 2304
rect 42524 2320 42576 2372
rect 56048 2388 56100 2440
rect 56416 2363 56468 2372
rect 56416 2329 56425 2363
rect 56425 2329 56459 2363
rect 56459 2329 56468 2363
rect 65064 2388 65116 2440
rect 56416 2320 56468 2329
rect 67640 2320 67692 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 26608 1980 26660 2032
rect 56416 1980 56468 2032
rect 50620 1300 50672 1352
rect 66168 1300 66220 1352
<< metal2 >>
rect 634 71200 746 72000
rect 1278 71200 1390 72000
rect 2566 71200 2678 72000
rect 3854 71346 3966 72000
rect 2976 71318 3966 71346
rect 1398 70952 1454 70961
rect 1398 70887 1454 70896
rect 1412 69426 1440 70887
rect 1400 69420 1452 69426
rect 1400 69362 1452 69368
rect 1584 69352 1636 69358
rect 1584 69294 1636 69300
rect 1596 67250 1624 69294
rect 2504 69216 2556 69222
rect 2504 69158 2556 69164
rect 2516 68882 2544 69158
rect 2504 68876 2556 68882
rect 2504 68818 2556 68824
rect 2780 68876 2832 68882
rect 2780 68818 2832 68824
rect 2792 68785 2820 68818
rect 2778 68776 2834 68785
rect 1860 68740 1912 68746
rect 2778 68711 2834 68720
rect 1860 68682 1912 68688
rect 1872 68474 1900 68682
rect 1860 68468 1912 68474
rect 1860 68410 1912 68416
rect 2044 68332 2096 68338
rect 2044 68274 2096 68280
rect 2056 67726 2084 68274
rect 2320 67788 2372 67794
rect 2320 67730 2372 67736
rect 2044 67720 2096 67726
rect 2044 67662 2096 67668
rect 2056 67250 2084 67662
rect 2332 67658 2360 67730
rect 2320 67652 2372 67658
rect 2320 67594 2372 67600
rect 1584 67244 1636 67250
rect 1584 67186 1636 67192
rect 2044 67244 2096 67250
rect 2044 67186 2096 67192
rect 1400 66632 1452 66638
rect 1400 66574 1452 66580
rect 1412 64666 1440 66574
rect 1584 66564 1636 66570
rect 1584 66506 1636 66512
rect 1596 66298 1624 66506
rect 1584 66292 1636 66298
rect 1584 66234 1636 66240
rect 1768 65544 1820 65550
rect 1768 65486 1820 65492
rect 1780 65074 1808 65486
rect 1952 65408 2004 65414
rect 1952 65350 2004 65356
rect 1964 65142 1992 65350
rect 1952 65136 2004 65142
rect 1952 65078 2004 65084
rect 1768 65068 1820 65074
rect 1768 65010 1820 65016
rect 1400 64660 1452 64666
rect 1400 64602 1452 64608
rect 1400 63368 1452 63374
rect 1398 63336 1400 63345
rect 1452 63336 1454 63345
rect 1398 63271 1454 63280
rect 1860 60784 1912 60790
rect 1860 60726 1912 60732
rect 1872 60625 1900 60726
rect 1858 60616 1914 60625
rect 1858 60551 1914 60560
rect 2136 60512 2188 60518
rect 2136 60454 2188 60460
rect 1676 60104 1728 60110
rect 1676 60046 1728 60052
rect 1688 59634 1716 60046
rect 1676 59628 1728 59634
rect 1676 59570 1728 59576
rect 1860 59560 1912 59566
rect 1860 59502 1912 59508
rect 1872 59226 1900 59502
rect 1860 59220 1912 59226
rect 1860 59162 1912 59168
rect 2044 59016 2096 59022
rect 2044 58958 2096 58964
rect 1400 56840 1452 56846
rect 1400 56782 1452 56788
rect 1412 56545 1440 56782
rect 1492 56704 1544 56710
rect 1492 56646 1544 56652
rect 1398 56536 1454 56545
rect 1398 56471 1454 56480
rect 1400 52896 1452 52902
rect 1400 52838 1452 52844
rect 1412 52562 1440 52838
rect 1400 52556 1452 52562
rect 1400 52498 1452 52504
rect 1504 45554 1532 56646
rect 1952 53984 2004 53990
rect 1952 53926 2004 53932
rect 1964 53650 1992 53926
rect 1952 53644 2004 53650
rect 1952 53586 2004 53592
rect 1860 52556 1912 52562
rect 1860 52498 1912 52504
rect 1872 52465 1900 52498
rect 1858 52456 1914 52465
rect 1584 52420 1636 52426
rect 1858 52391 1914 52400
rect 1584 52362 1636 52368
rect 1596 52154 1624 52362
rect 1584 52148 1636 52154
rect 1584 52090 1636 52096
rect 2056 52018 2084 58958
rect 2148 56506 2176 60454
rect 2136 56500 2188 56506
rect 2136 56442 2188 56448
rect 2044 52012 2096 52018
rect 2044 51954 2096 51960
rect 1676 48136 1728 48142
rect 1676 48078 1728 48084
rect 1688 47666 1716 48078
rect 1676 47660 1728 47666
rect 1676 47602 1728 47608
rect 2332 47054 2360 67594
rect 2778 67416 2834 67425
rect 2778 67351 2834 67360
rect 2596 67244 2648 67250
rect 2596 67186 2648 67192
rect 2608 66162 2636 67186
rect 2792 66706 2820 67351
rect 2872 67176 2924 67182
rect 2872 67118 2924 67124
rect 2780 66700 2832 66706
rect 2780 66642 2832 66648
rect 2596 66156 2648 66162
rect 2596 66098 2648 66104
rect 2884 65482 2912 67118
rect 2872 65476 2924 65482
rect 2872 65418 2924 65424
rect 2976 61878 3004 71318
rect 3854 71200 3966 71318
rect 5142 71200 5254 72000
rect 6430 71200 6542 72000
rect 7718 71200 7830 72000
rect 9006 71200 9118 72000
rect 10294 71200 10406 72000
rect 11582 71200 11694 72000
rect 12870 71200 12982 72000
rect 14158 71200 14270 72000
rect 15446 71200 15558 72000
rect 16734 71200 16846 72000
rect 18022 71200 18134 72000
rect 19310 71200 19422 72000
rect 20598 71200 20710 72000
rect 21886 71200 21998 72000
rect 23174 71346 23286 72000
rect 22112 71318 23286 71346
rect 4804 69216 4856 69222
rect 4804 69158 4856 69164
rect 4214 69116 4522 69136
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69040 4522 69060
rect 4620 68808 4672 68814
rect 4620 68750 4672 68756
rect 4632 68474 4660 68750
rect 4712 68672 4764 68678
rect 4712 68614 4764 68620
rect 4620 68468 4672 68474
rect 4620 68410 4672 68416
rect 3056 68264 3108 68270
rect 3056 68206 3108 68212
rect 3332 68264 3384 68270
rect 3332 68206 3384 68212
rect 3068 67182 3096 68206
rect 3056 67176 3108 67182
rect 3056 67118 3108 67124
rect 3068 64874 3096 67118
rect 3068 64846 3188 64874
rect 2964 61872 3016 61878
rect 2964 61814 3016 61820
rect 2780 59560 2832 59566
rect 2780 59502 2832 59508
rect 2792 59265 2820 59502
rect 2778 59256 2834 59265
rect 2778 59191 2834 59200
rect 2778 53816 2834 53825
rect 2778 53751 2834 53760
rect 2792 53650 2820 53751
rect 2780 53644 2832 53650
rect 2780 53586 2832 53592
rect 2412 53508 2464 53514
rect 2412 53450 2464 53456
rect 2424 53242 2452 53450
rect 2412 53236 2464 53242
rect 2412 53178 2464 53184
rect 2778 47696 2834 47705
rect 2778 47631 2834 47640
rect 2792 47598 2820 47631
rect 2412 47592 2464 47598
rect 2412 47534 2464 47540
rect 2780 47592 2832 47598
rect 2780 47534 2832 47540
rect 2424 47258 2452 47534
rect 2412 47252 2464 47258
rect 2412 47194 2464 47200
rect 2320 47048 2372 47054
rect 2320 46990 2372 46996
rect 1860 46572 1912 46578
rect 1860 46514 1912 46520
rect 1872 46345 1900 46514
rect 2044 46436 2096 46442
rect 2044 46378 2096 46384
rect 1858 46336 1914 46345
rect 1858 46271 1914 46280
rect 1504 45526 1716 45554
rect 1400 39840 1452 39846
rect 1400 39782 1452 39788
rect 1412 39506 1440 39782
rect 1400 39500 1452 39506
rect 1400 39442 1452 39448
rect 20 37732 72 37738
rect 20 37674 72 37680
rect 32 800 60 37674
rect 1584 36576 1636 36582
rect 1584 36518 1636 36524
rect 1596 36242 1624 36518
rect 1584 36236 1636 36242
rect 1584 36178 1636 36184
rect 1400 36168 1452 36174
rect 1400 36110 1452 36116
rect 1412 35698 1440 36110
rect 1400 35692 1452 35698
rect 1400 35634 1452 35640
rect 1688 35494 1716 45526
rect 1860 45484 1912 45490
rect 1860 45426 1912 45432
rect 1872 44985 1900 45426
rect 1952 45280 2004 45286
rect 1952 45222 2004 45228
rect 1964 45082 1992 45222
rect 1952 45076 2004 45082
rect 1952 45018 2004 45024
rect 1858 44976 1914 44985
rect 1858 44911 1914 44920
rect 1860 43716 1912 43722
rect 1860 43658 1912 43664
rect 1872 43625 1900 43658
rect 1858 43616 1914 43625
rect 1858 43551 1914 43560
rect 1860 42628 1912 42634
rect 1860 42570 1912 42576
rect 1872 42265 1900 42570
rect 1952 42560 2004 42566
rect 1952 42502 2004 42508
rect 1964 42362 1992 42502
rect 1952 42356 2004 42362
rect 1952 42298 2004 42304
rect 2056 42265 2084 46378
rect 1858 42256 1914 42265
rect 1858 42191 1914 42200
rect 2042 42256 2098 42265
rect 2042 42191 2098 42200
rect 2778 39536 2834 39545
rect 2778 39471 2780 39480
rect 2832 39471 2834 39480
rect 2780 39442 2832 39448
rect 1860 39364 1912 39370
rect 1860 39306 1912 39312
rect 1872 39098 1900 39306
rect 1860 39092 1912 39098
rect 1860 39034 1912 39040
rect 3160 38962 3188 64846
rect 3238 40896 3294 40905
rect 3238 40831 3294 40840
rect 3252 40458 3280 40831
rect 3240 40452 3292 40458
rect 3240 40394 3292 40400
rect 3148 38956 3200 38962
rect 3148 38898 3200 38904
rect 3240 38548 3292 38554
rect 3240 38490 3292 38496
rect 3252 38185 3280 38490
rect 3238 38176 3294 38185
rect 3238 38111 3294 38120
rect 3240 37188 3292 37194
rect 3240 37130 3292 37136
rect 3252 36825 3280 37130
rect 3238 36816 3294 36825
rect 3238 36751 3294 36760
rect 2780 36236 2832 36242
rect 2780 36178 2832 36184
rect 1676 35488 1728 35494
rect 2792 35465 2820 36178
rect 1676 35430 1728 35436
rect 2778 35456 2834 35465
rect 2778 35391 2834 35400
rect 1400 34536 1452 34542
rect 1400 34478 1452 34484
rect 1412 34105 1440 34478
rect 1398 34096 1454 34105
rect 1398 34031 1454 34040
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 1688 31346 1716 31758
rect 2778 31376 2834 31385
rect 1676 31340 1728 31346
rect 2778 31311 2834 31320
rect 1676 31282 1728 31288
rect 2792 31278 2820 31311
rect 2044 31272 2096 31278
rect 2044 31214 2096 31220
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2056 30938 2084 31214
rect 2044 30932 2096 30938
rect 2044 30874 2096 30880
rect 3344 30734 3372 68206
rect 4214 68028 4522 68048
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67952 4522 67972
rect 4214 66940 4522 66960
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66864 4522 66884
rect 4068 66632 4120 66638
rect 4068 66574 4120 66580
rect 4080 66162 4108 66574
rect 4068 66156 4120 66162
rect 4068 66098 4120 66104
rect 3424 66020 3476 66026
rect 3424 65962 3476 65968
rect 1952 30728 2004 30734
rect 1952 30670 2004 30676
rect 3332 30728 3384 30734
rect 3332 30670 3384 30676
rect 1860 30184 1912 30190
rect 1860 30126 1912 30132
rect 1872 29850 1900 30126
rect 1860 29844 1912 29850
rect 1860 29786 1912 29792
rect 1676 26376 1728 26382
rect 1676 26318 1728 26324
rect 1688 25906 1716 26318
rect 1676 25900 1728 25906
rect 1676 25842 1728 25848
rect 1860 24812 1912 24818
rect 1860 24754 1912 24760
rect 1872 24585 1900 24754
rect 1858 24576 1914 24585
rect 1858 24511 1914 24520
rect 1768 22568 1820 22574
rect 1768 22510 1820 22516
rect 1780 22234 1808 22510
rect 1768 22228 1820 22234
rect 1768 22170 1820 22176
rect 1860 21548 1912 21554
rect 1860 21490 1912 21496
rect 1872 21185 1900 21490
rect 1858 21176 1914 21185
rect 1858 21111 1914 21120
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1596 12850 1624 13262
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1780 12442 1808 12718
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1872 7585 1900 7754
rect 1858 7576 1914 7585
rect 1858 7511 1914 7520
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 664 3732 716 3738
rect 664 3674 716 3680
rect 676 800 704 3674
rect 1596 3058 1624 3878
rect 1964 3534 1992 30670
rect 2780 30184 2832 30190
rect 2780 30126 2832 30132
rect 2872 30184 2924 30190
rect 2872 30126 2924 30132
rect 2792 29850 2820 30126
rect 2884 30025 2912 30126
rect 2870 30016 2926 30025
rect 2870 29951 2926 29960
rect 2780 29844 2832 29850
rect 2780 29786 2832 29792
rect 3054 27296 3110 27305
rect 3054 27231 3110 27240
rect 3068 26382 3096 27231
rect 3056 26376 3108 26382
rect 3056 26318 3108 26324
rect 2778 25936 2834 25945
rect 2778 25871 2834 25880
rect 2792 25838 2820 25871
rect 2320 25832 2372 25838
rect 2320 25774 2372 25780
rect 2780 25832 2832 25838
rect 2780 25774 2832 25780
rect 2332 25498 2360 25774
rect 2320 25492 2372 25498
rect 2320 25434 2372 25440
rect 3436 25294 3464 65962
rect 4080 65550 4108 66098
rect 4214 65852 4522 65872
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65776 4522 65796
rect 4068 65544 4120 65550
rect 4068 65486 4120 65492
rect 4080 65074 4108 65486
rect 4344 65476 4396 65482
rect 4344 65418 4396 65424
rect 4068 65068 4120 65074
rect 4068 65010 4120 65016
rect 4356 65006 4384 65418
rect 3608 65000 3660 65006
rect 3608 64942 3660 64948
rect 4344 65000 4396 65006
rect 4344 64942 4396 64948
rect 3514 55176 3570 55185
rect 3514 55111 3570 55120
rect 3528 54058 3556 55111
rect 3516 54052 3568 54058
rect 3516 53994 3568 54000
rect 3516 52420 3568 52426
rect 3516 52362 3568 52368
rect 3528 51105 3556 52362
rect 3514 51096 3570 51105
rect 3514 51031 3570 51040
rect 3516 49972 3568 49978
rect 3516 49914 3568 49920
rect 3528 49745 3556 49914
rect 3514 49736 3570 49745
rect 3514 49671 3570 49680
rect 3424 25288 3476 25294
rect 3424 25230 3476 25236
rect 2044 24608 2096 24614
rect 2044 24550 2096 24556
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 2056 24274 2084 24550
rect 3436 24342 3464 24550
rect 3424 24336 3476 24342
rect 3424 24278 3476 24284
rect 2044 24268 2096 24274
rect 2044 24210 2096 24216
rect 2780 24268 2832 24274
rect 2780 24210 2832 24216
rect 2792 23905 2820 24210
rect 2778 23896 2834 23905
rect 2778 23831 2834 23840
rect 2596 22568 2648 22574
rect 2780 22568 2832 22574
rect 2596 22510 2648 22516
rect 2778 22536 2780 22545
rect 2832 22536 2834 22545
rect 2608 22234 2636 22510
rect 2778 22471 2834 22480
rect 2596 22228 2648 22234
rect 2596 22170 2648 22176
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2964 16040 3016 16046
rect 2964 15982 3016 15988
rect 2056 15706 2084 15982
rect 2884 15706 2912 15982
rect 2976 15745 3004 15982
rect 2962 15736 3018 15745
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2872 15700 2924 15706
rect 2962 15671 3018 15680
rect 2872 15642 2924 15648
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2778 13016 2834 13025
rect 2778 12951 2834 12960
rect 2792 12782 2820 12951
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1780 3126 1808 3334
rect 1964 3194 1992 3470
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 1768 3120 1820 3126
rect 1768 3062 1820 3068
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 2424 2446 2452 12174
rect 2884 6914 2912 15438
rect 2792 6886 2912 6914
rect 2792 5710 2820 6886
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 3620 4865 3648 64942
rect 4214 64764 4522 64784
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64688 4522 64708
rect 4214 63676 4522 63696
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63600 4522 63620
rect 4214 62588 4522 62608
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62512 4522 62532
rect 4214 61500 4522 61520
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61424 4522 61444
rect 4214 60412 4522 60432
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60336 4522 60356
rect 4214 59324 4522 59344
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59248 4522 59268
rect 4214 58236 4522 58256
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58160 4522 58180
rect 4214 57148 4522 57168
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57072 4522 57092
rect 4214 56060 4522 56080
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55984 4522 56004
rect 4214 54972 4522 54992
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54896 4522 54916
rect 4214 53884 4522 53904
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53808 4522 53828
rect 4214 52796 4522 52816
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52720 4522 52740
rect 4214 51708 4522 51728
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51632 4522 51652
rect 4214 50620 4522 50640
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50544 4522 50564
rect 4214 49532 4522 49552
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49456 4522 49476
rect 4214 48444 4522 48464
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48368 4522 48388
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4632 22030 4660 68410
rect 4724 67794 4752 68614
rect 4816 67862 4844 69158
rect 4804 67856 4856 67862
rect 4804 67798 4856 67804
rect 5184 67794 5212 71200
rect 6000 69216 6052 69222
rect 6000 69158 6052 69164
rect 6012 68882 6040 69158
rect 6472 68882 6500 71200
rect 7760 69426 7788 71200
rect 7748 69420 7800 69426
rect 7748 69362 7800 69368
rect 8024 69216 8076 69222
rect 8024 69158 8076 69164
rect 6000 68876 6052 68882
rect 6000 68818 6052 68824
rect 6460 68876 6512 68882
rect 6460 68818 6512 68824
rect 5908 68808 5960 68814
rect 5908 68750 5960 68756
rect 4712 67788 4764 67794
rect 4712 67730 4764 67736
rect 5172 67788 5224 67794
rect 5172 67730 5224 67736
rect 5172 67176 5224 67182
rect 5172 67118 5224 67124
rect 4712 66496 4764 66502
rect 4712 66438 4764 66444
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 3976 18148 4028 18154
rect 3976 18090 4028 18096
rect 3606 4856 3662 4865
rect 3606 4791 3662 4800
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3160 3505 3188 3606
rect 3884 3528 3936 3534
rect 3146 3496 3202 3505
rect 3884 3470 3936 3476
rect 3146 3431 3202 3440
rect 3896 3058 3924 3470
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 2792 2145 2820 2926
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect -10 0 102 800
rect 634 0 746 800
rect 1922 0 2034 800
rect 2884 785 2912 2858
rect 3528 2650 3556 2926
rect 3988 2650 4016 18090
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4724 15502 4752 66438
rect 4804 65476 4856 65482
rect 4804 65418 4856 65424
rect 4816 65210 4844 65418
rect 4804 65204 4856 65210
rect 4804 65146 4856 65152
rect 4816 29646 4844 65146
rect 5184 53106 5212 67118
rect 5920 66706 5948 68750
rect 5908 66700 5960 66706
rect 5908 66642 5960 66648
rect 5264 66088 5316 66094
rect 5264 66030 5316 66036
rect 5172 53100 5224 53106
rect 5172 53042 5224 53048
rect 4804 29640 4856 29646
rect 4804 29582 4856 29588
rect 5276 24818 5304 66030
rect 5920 64874 5948 66642
rect 5920 64846 6040 64874
rect 6012 59022 6040 64846
rect 6000 59016 6052 59022
rect 6000 58958 6052 58964
rect 6552 54120 6604 54126
rect 6552 54062 6604 54068
rect 6564 53786 6592 54062
rect 6552 53780 6604 53786
rect 6552 53722 6604 53728
rect 6368 53576 6420 53582
rect 6368 53518 6420 53524
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 6380 4690 6408 53518
rect 6828 47048 6880 47054
rect 6828 46990 6880 46996
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6380 4554 6408 4626
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6380 4146 6408 4490
rect 6840 4146 6868 46990
rect 8036 35562 8064 69158
rect 11624 68950 11652 71200
rect 14200 69494 14228 71200
rect 14188 69488 14240 69494
rect 14188 69430 14240 69436
rect 14832 69284 14884 69290
rect 14832 69226 14884 69232
rect 11704 69216 11756 69222
rect 11704 69158 11756 69164
rect 11612 68944 11664 68950
rect 11612 68886 11664 68892
rect 11716 68882 11744 69158
rect 11704 68876 11756 68882
rect 11704 68818 11756 68824
rect 10416 68808 10468 68814
rect 10416 68750 10468 68756
rect 10428 66706 10456 68750
rect 10416 66700 10468 66706
rect 10416 66642 10468 66648
rect 14648 59628 14700 59634
rect 14648 59570 14700 59576
rect 14372 59424 14424 59430
rect 14372 59366 14424 59372
rect 14384 59022 14412 59366
rect 14096 59016 14148 59022
rect 14096 58958 14148 58964
rect 14372 59016 14424 59022
rect 14372 58958 14424 58964
rect 14108 58682 14136 58958
rect 14660 58682 14688 59570
rect 14096 58676 14148 58682
rect 14096 58618 14148 58624
rect 14648 58676 14700 58682
rect 14648 58618 14700 58624
rect 13820 58540 13872 58546
rect 13820 58482 13872 58488
rect 13832 56846 13860 58482
rect 14372 57384 14424 57390
rect 14372 57326 14424 57332
rect 14384 57050 14412 57326
rect 14372 57044 14424 57050
rect 14372 56986 14424 56992
rect 13820 56840 13872 56846
rect 13820 56782 13872 56788
rect 13832 55282 13860 56782
rect 14648 55616 14700 55622
rect 14648 55558 14700 55564
rect 14660 55350 14688 55558
rect 14648 55344 14700 55350
rect 14648 55286 14700 55292
rect 13820 55276 13872 55282
rect 13820 55218 13872 55224
rect 13832 53582 13860 55218
rect 13820 53576 13872 53582
rect 13820 53518 13872 53524
rect 13544 53440 13596 53446
rect 13544 53382 13596 53388
rect 13556 53106 13584 53382
rect 13544 53100 13596 53106
rect 13544 53042 13596 53048
rect 13832 51270 13860 53518
rect 14280 53440 14332 53446
rect 14280 53382 14332 53388
rect 14096 53100 14148 53106
rect 14096 53042 14148 53048
rect 14108 52698 14136 53042
rect 14096 52692 14148 52698
rect 14096 52634 14148 52640
rect 14292 52494 14320 53382
rect 14280 52488 14332 52494
rect 14280 52430 14332 52436
rect 14372 51944 14424 51950
rect 14372 51886 14424 51892
rect 13820 51264 13872 51270
rect 13820 51206 13872 51212
rect 14384 51066 14412 51886
rect 14648 51264 14700 51270
rect 14648 51206 14700 51212
rect 14740 51264 14792 51270
rect 14740 51206 14792 51212
rect 14372 51060 14424 51066
rect 14372 51002 14424 51008
rect 14660 50930 14688 51206
rect 14096 50924 14148 50930
rect 14096 50866 14148 50872
rect 14648 50924 14700 50930
rect 14648 50866 14700 50872
rect 14108 50318 14136 50866
rect 14280 50720 14332 50726
rect 14280 50662 14332 50668
rect 14096 50312 14148 50318
rect 14096 50254 14148 50260
rect 13820 50244 13872 50250
rect 13820 50186 13872 50192
rect 12440 50176 12492 50182
rect 12440 50118 12492 50124
rect 12452 49842 12480 50118
rect 12440 49836 12492 49842
rect 12440 49778 12492 49784
rect 12992 49836 13044 49842
rect 12992 49778 13044 49784
rect 13004 48890 13032 49778
rect 13832 49706 13860 50186
rect 13820 49700 13872 49706
rect 13820 49642 13872 49648
rect 13832 49298 13860 49642
rect 13820 49292 13872 49298
rect 13820 49234 13872 49240
rect 13268 49224 13320 49230
rect 13268 49166 13320 49172
rect 13176 49088 13228 49094
rect 13176 49030 13228 49036
rect 12992 48884 13044 48890
rect 12992 48826 13044 48832
rect 13188 48754 13216 49030
rect 13280 48822 13308 49166
rect 13268 48816 13320 48822
rect 13268 48758 13320 48764
rect 13176 48748 13228 48754
rect 13176 48690 13228 48696
rect 12716 48000 12768 48006
rect 12716 47942 12768 47948
rect 12728 47734 12756 47942
rect 12716 47728 12768 47734
rect 12716 47670 12768 47676
rect 12164 47592 12216 47598
rect 12164 47534 12216 47540
rect 12176 47258 12204 47534
rect 12164 47252 12216 47258
rect 12164 47194 12216 47200
rect 13280 47054 13308 48758
rect 14108 48550 14136 50254
rect 14292 49842 14320 50662
rect 14280 49836 14332 49842
rect 14280 49778 14332 49784
rect 14372 49836 14424 49842
rect 14372 49778 14424 49784
rect 14384 49434 14412 49778
rect 14372 49428 14424 49434
rect 14372 49370 14424 49376
rect 14096 48544 14148 48550
rect 14096 48486 14148 48492
rect 13360 48136 13412 48142
rect 13360 48078 13412 48084
rect 13372 47258 13400 48078
rect 13544 47456 13596 47462
rect 13544 47398 13596 47404
rect 13360 47252 13412 47258
rect 13360 47194 13412 47200
rect 13556 47122 13584 47398
rect 14108 47190 14136 48486
rect 14464 48136 14516 48142
rect 14464 48078 14516 48084
rect 14188 48000 14240 48006
rect 14188 47942 14240 47948
rect 14200 47666 14228 47942
rect 14188 47660 14240 47666
rect 14188 47602 14240 47608
rect 14096 47184 14148 47190
rect 14096 47126 14148 47132
rect 13544 47116 13596 47122
rect 13544 47058 13596 47064
rect 12624 47048 12676 47054
rect 12624 46990 12676 46996
rect 13268 47048 13320 47054
rect 13268 46990 13320 46996
rect 12532 45416 12584 45422
rect 12532 45358 12584 45364
rect 12544 45082 12572 45358
rect 12532 45076 12584 45082
rect 12532 45018 12584 45024
rect 12636 44878 12664 46990
rect 12992 45824 13044 45830
rect 12992 45766 13044 45772
rect 13004 45558 13032 45766
rect 12992 45552 13044 45558
rect 13280 45554 13308 46990
rect 14476 45966 14504 48078
rect 13544 45960 13596 45966
rect 13544 45902 13596 45908
rect 14464 45960 14516 45966
rect 14464 45902 14516 45908
rect 13280 45526 13400 45554
rect 12992 45494 13044 45500
rect 13176 45280 13228 45286
rect 13176 45222 13228 45228
rect 13188 44946 13216 45222
rect 13176 44940 13228 44946
rect 13176 44882 13228 44888
rect 13372 44878 13400 45526
rect 13556 45082 13584 45902
rect 14476 45554 14504 45902
rect 14648 45824 14700 45830
rect 14648 45766 14700 45772
rect 14476 45526 14596 45554
rect 13544 45076 13596 45082
rect 13544 45018 13596 45024
rect 12624 44872 12676 44878
rect 12624 44814 12676 44820
rect 13360 44872 13412 44878
rect 13360 44814 13412 44820
rect 12636 44402 12664 44814
rect 12624 44396 12676 44402
rect 12624 44338 12676 44344
rect 12624 44192 12676 44198
rect 12624 44134 12676 44140
rect 12636 43314 12664 44134
rect 13372 43790 13400 44814
rect 14568 44538 14596 45526
rect 14660 45490 14688 45766
rect 14648 45484 14700 45490
rect 14648 45426 14700 45432
rect 14556 44532 14608 44538
rect 14556 44474 14608 44480
rect 13360 43784 13412 43790
rect 13360 43726 13412 43732
rect 14096 43716 14148 43722
rect 14096 43658 14148 43664
rect 13360 43648 13412 43654
rect 13360 43590 13412 43596
rect 12624 43308 12676 43314
rect 12624 43250 12676 43256
rect 12992 43308 13044 43314
rect 12992 43250 13044 43256
rect 13004 42906 13032 43250
rect 12992 42900 13044 42906
rect 12992 42842 13044 42848
rect 13372 42702 13400 43590
rect 14108 43178 14136 43658
rect 14568 43314 14596 44474
rect 14752 44402 14780 51206
rect 14740 44396 14792 44402
rect 14740 44338 14792 44344
rect 14648 43784 14700 43790
rect 14648 43726 14700 43732
rect 14660 43450 14688 43726
rect 14648 43444 14700 43450
rect 14648 43386 14700 43392
rect 14556 43308 14608 43314
rect 14556 43250 14608 43256
rect 14096 43172 14148 43178
rect 14096 43114 14148 43120
rect 14568 42702 14596 43250
rect 13360 42696 13412 42702
rect 13360 42638 13412 42644
rect 14556 42696 14608 42702
rect 14556 42638 14608 42644
rect 14740 42560 14792 42566
rect 14740 42502 14792 42508
rect 14752 42226 14780 42502
rect 14740 42220 14792 42226
rect 14740 42162 14792 42168
rect 14844 41750 14872 69226
rect 16776 68950 16804 71200
rect 19352 69494 19380 71200
rect 19574 69660 19882 69680
rect 19574 69658 19580 69660
rect 19636 69658 19660 69660
rect 19716 69658 19740 69660
rect 19796 69658 19820 69660
rect 19876 69658 19882 69660
rect 19636 69606 19638 69658
rect 19818 69606 19820 69658
rect 19574 69604 19580 69606
rect 19636 69604 19660 69606
rect 19716 69604 19740 69606
rect 19796 69604 19820 69606
rect 19876 69604 19882 69606
rect 19574 69584 19882 69604
rect 20640 69494 20668 71200
rect 19340 69488 19392 69494
rect 19340 69430 19392 69436
rect 20628 69488 20680 69494
rect 20628 69430 20680 69436
rect 20260 69284 20312 69290
rect 20260 69226 20312 69232
rect 21640 69284 21692 69290
rect 21640 69226 21692 69232
rect 16856 69216 16908 69222
rect 16856 69158 16908 69164
rect 16764 68944 16816 68950
rect 16764 68886 16816 68892
rect 16868 68882 16896 69158
rect 16856 68876 16908 68882
rect 16856 68818 16908 68824
rect 15476 68808 15528 68814
rect 15476 68750 15528 68756
rect 15488 68678 15516 68750
rect 15476 68672 15528 68678
rect 15476 68614 15528 68620
rect 15488 65006 15516 68614
rect 19574 68572 19882 68592
rect 19574 68570 19580 68572
rect 19636 68570 19660 68572
rect 19716 68570 19740 68572
rect 19796 68570 19820 68572
rect 19876 68570 19882 68572
rect 19636 68518 19638 68570
rect 19818 68518 19820 68570
rect 19574 68516 19580 68518
rect 19636 68516 19660 68518
rect 19716 68516 19740 68518
rect 19796 68516 19820 68518
rect 19876 68516 19882 68518
rect 19574 68496 19882 68516
rect 19574 67484 19882 67504
rect 19574 67482 19580 67484
rect 19636 67482 19660 67484
rect 19716 67482 19740 67484
rect 19796 67482 19820 67484
rect 19876 67482 19882 67484
rect 19636 67430 19638 67482
rect 19818 67430 19820 67482
rect 19574 67428 19580 67430
rect 19636 67428 19660 67430
rect 19716 67428 19740 67430
rect 19796 67428 19820 67430
rect 19876 67428 19882 67430
rect 19574 67408 19882 67428
rect 19574 66396 19882 66416
rect 19574 66394 19580 66396
rect 19636 66394 19660 66396
rect 19716 66394 19740 66396
rect 19796 66394 19820 66396
rect 19876 66394 19882 66396
rect 19636 66342 19638 66394
rect 19818 66342 19820 66394
rect 19574 66340 19580 66342
rect 19636 66340 19660 66342
rect 19716 66340 19740 66342
rect 19796 66340 19820 66342
rect 19876 66340 19882 66342
rect 19574 66320 19882 66340
rect 19574 65308 19882 65328
rect 19574 65306 19580 65308
rect 19636 65306 19660 65308
rect 19716 65306 19740 65308
rect 19796 65306 19820 65308
rect 19876 65306 19882 65308
rect 19636 65254 19638 65306
rect 19818 65254 19820 65306
rect 19574 65252 19580 65254
rect 19636 65252 19660 65254
rect 19716 65252 19740 65254
rect 19796 65252 19820 65254
rect 19876 65252 19882 65254
rect 19574 65232 19882 65252
rect 15476 65000 15528 65006
rect 15476 64942 15528 64948
rect 19574 64220 19882 64240
rect 19574 64218 19580 64220
rect 19636 64218 19660 64220
rect 19716 64218 19740 64220
rect 19796 64218 19820 64220
rect 19876 64218 19882 64220
rect 19636 64166 19638 64218
rect 19818 64166 19820 64218
rect 19574 64164 19580 64166
rect 19636 64164 19660 64166
rect 19716 64164 19740 64166
rect 19796 64164 19820 64166
rect 19876 64164 19882 64166
rect 19574 64144 19882 64164
rect 19574 63132 19882 63152
rect 19574 63130 19580 63132
rect 19636 63130 19660 63132
rect 19716 63130 19740 63132
rect 19796 63130 19820 63132
rect 19876 63130 19882 63132
rect 19636 63078 19638 63130
rect 19818 63078 19820 63130
rect 19574 63076 19580 63078
rect 19636 63076 19660 63078
rect 19716 63076 19740 63078
rect 19796 63076 19820 63078
rect 19876 63076 19882 63078
rect 19574 63056 19882 63076
rect 19340 62144 19392 62150
rect 19340 62086 19392 62092
rect 19352 61946 19380 62086
rect 19574 62044 19882 62064
rect 19574 62042 19580 62044
rect 19636 62042 19660 62044
rect 19716 62042 19740 62044
rect 19796 62042 19820 62044
rect 19876 62042 19882 62044
rect 19636 61990 19638 62042
rect 19818 61990 19820 62042
rect 19574 61988 19580 61990
rect 19636 61988 19660 61990
rect 19716 61988 19740 61990
rect 19796 61988 19820 61990
rect 19876 61988 19882 61990
rect 19574 61968 19882 61988
rect 19340 61940 19392 61946
rect 19340 61882 19392 61888
rect 19340 61804 19392 61810
rect 19340 61746 19392 61752
rect 18236 61192 18288 61198
rect 18236 61134 18288 61140
rect 17040 60716 17092 60722
rect 17040 60658 17092 60664
rect 17500 60716 17552 60722
rect 17500 60658 17552 60664
rect 15844 60512 15896 60518
rect 15844 60454 15896 60460
rect 16028 60512 16080 60518
rect 16028 60454 16080 60460
rect 15856 60110 15884 60454
rect 15568 60104 15620 60110
rect 15568 60046 15620 60052
rect 15844 60104 15896 60110
rect 15844 60046 15896 60052
rect 15580 59770 15608 60046
rect 15568 59764 15620 59770
rect 15568 59706 15620 59712
rect 15844 59628 15896 59634
rect 15844 59570 15896 59576
rect 15476 59152 15528 59158
rect 15476 59094 15528 59100
rect 15488 58614 15516 59094
rect 15476 58608 15528 58614
rect 15476 58550 15528 58556
rect 15200 58540 15252 58546
rect 15200 58482 15252 58488
rect 14924 57452 14976 57458
rect 14924 57394 14976 57400
rect 14936 56234 14964 57394
rect 15212 56846 15240 58482
rect 15856 57934 15884 59570
rect 16040 58546 16068 60454
rect 16580 60104 16632 60110
rect 16580 60046 16632 60052
rect 16592 59634 16620 60046
rect 16948 59968 17000 59974
rect 16948 59910 17000 59916
rect 16580 59628 16632 59634
rect 16580 59570 16632 59576
rect 16028 58540 16080 58546
rect 16028 58482 16080 58488
rect 15844 57928 15896 57934
rect 15844 57870 15896 57876
rect 15752 57316 15804 57322
rect 15752 57258 15804 57264
rect 15764 56914 15792 57258
rect 15752 56908 15804 56914
rect 15752 56850 15804 56856
rect 15200 56840 15252 56846
rect 15200 56782 15252 56788
rect 14924 56228 14976 56234
rect 14924 56170 14976 56176
rect 15212 54670 15240 56782
rect 15384 56704 15436 56710
rect 15384 56646 15436 56652
rect 15396 56370 15424 56646
rect 15384 56364 15436 56370
rect 15384 56306 15436 56312
rect 15292 55752 15344 55758
rect 15292 55694 15344 55700
rect 15304 54874 15332 55694
rect 15568 55072 15620 55078
rect 15568 55014 15620 55020
rect 15292 54868 15344 54874
rect 15292 54810 15344 54816
rect 15200 54664 15252 54670
rect 15200 54606 15252 54612
rect 15212 53666 15240 54606
rect 15580 54602 15608 55014
rect 15568 54596 15620 54602
rect 15568 54538 15620 54544
rect 15212 53650 15332 53666
rect 15200 53644 15332 53650
rect 15252 53638 15332 53644
rect 15200 53586 15252 53592
rect 15200 53508 15252 53514
rect 15200 53450 15252 53456
rect 15212 52902 15240 53450
rect 15200 52896 15252 52902
rect 15200 52838 15252 52844
rect 15304 52698 15332 53638
rect 15568 53576 15620 53582
rect 15568 53518 15620 53524
rect 15580 53242 15608 53518
rect 15568 53236 15620 53242
rect 15568 53178 15620 53184
rect 15856 53106 15884 57870
rect 16592 57390 16620 59570
rect 16960 59566 16988 59910
rect 17052 59770 17080 60658
rect 17408 60648 17460 60654
rect 17408 60590 17460 60596
rect 17420 59770 17448 60590
rect 17040 59764 17092 59770
rect 17040 59706 17092 59712
rect 17408 59764 17460 59770
rect 17408 59706 17460 59712
rect 16948 59560 17000 59566
rect 16948 59502 17000 59508
rect 17512 59226 17540 60658
rect 17592 59968 17644 59974
rect 17592 59910 17644 59916
rect 17868 59968 17920 59974
rect 17868 59910 17920 59916
rect 17500 59220 17552 59226
rect 17500 59162 17552 59168
rect 17604 59022 17632 59910
rect 17880 59634 17908 59910
rect 17868 59628 17920 59634
rect 17868 59570 17920 59576
rect 17592 59016 17644 59022
rect 17592 58958 17644 58964
rect 17132 58540 17184 58546
rect 17132 58482 17184 58488
rect 16764 58336 16816 58342
rect 16764 58278 16816 58284
rect 16776 57934 16804 58278
rect 16764 57928 16816 57934
rect 16764 57870 16816 57876
rect 17144 57594 17172 58482
rect 17868 57792 17920 57798
rect 17868 57734 17920 57740
rect 17132 57588 17184 57594
rect 17132 57530 17184 57536
rect 17880 57526 17908 57734
rect 17868 57520 17920 57526
rect 17868 57462 17920 57468
rect 16580 57384 16632 57390
rect 16580 57326 16632 57332
rect 18144 57384 18196 57390
rect 18144 57326 18196 57332
rect 16028 56296 16080 56302
rect 16028 56238 16080 56244
rect 16040 55962 16068 56238
rect 16028 55956 16080 55962
rect 16028 55898 16080 55904
rect 16592 54194 16620 57326
rect 17960 57248 18012 57254
rect 17960 57190 18012 57196
rect 16948 56704 17000 56710
rect 16948 56646 17000 56652
rect 16960 56438 16988 56646
rect 16948 56432 17000 56438
rect 16948 56374 17000 56380
rect 17316 55752 17368 55758
rect 17316 55694 17368 55700
rect 16948 55616 17000 55622
rect 16948 55558 17000 55564
rect 16960 55282 16988 55558
rect 16948 55276 17000 55282
rect 16948 55218 17000 55224
rect 16580 54188 16632 54194
rect 16580 54130 16632 54136
rect 15844 53100 15896 53106
rect 15844 53042 15896 53048
rect 16304 52896 16356 52902
rect 16304 52838 16356 52844
rect 15292 52692 15344 52698
rect 15292 52634 15344 52640
rect 16316 52426 16344 52838
rect 16592 52562 16620 54130
rect 16856 53984 16908 53990
rect 16856 53926 16908 53932
rect 16948 53984 17000 53990
rect 16948 53926 17000 53932
rect 16672 53508 16724 53514
rect 16672 53450 16724 53456
rect 16684 53242 16712 53450
rect 16672 53236 16724 53242
rect 16672 53178 16724 53184
rect 16764 53168 16816 53174
rect 16764 53110 16816 53116
rect 16580 52556 16632 52562
rect 16580 52498 16632 52504
rect 16028 52420 16080 52426
rect 16028 52362 16080 52368
rect 16304 52420 16356 52426
rect 16304 52362 16356 52368
rect 15016 52012 15068 52018
rect 15016 51954 15068 51960
rect 15028 51610 15056 51954
rect 15752 51808 15804 51814
rect 15752 51750 15804 51756
rect 15016 51604 15068 51610
rect 15016 51546 15068 51552
rect 15764 51406 15792 51750
rect 15752 51400 15804 51406
rect 15752 51342 15804 51348
rect 15108 50312 15160 50318
rect 15108 50254 15160 50260
rect 15200 50312 15252 50318
rect 15200 50254 15252 50260
rect 15120 49842 15148 50254
rect 15108 49836 15160 49842
rect 15108 49778 15160 49784
rect 15212 49230 15240 50254
rect 15384 50176 15436 50182
rect 15384 50118 15436 50124
rect 15396 49298 15424 50118
rect 15384 49292 15436 49298
rect 15384 49234 15436 49240
rect 15200 49224 15252 49230
rect 15200 49166 15252 49172
rect 15016 48000 15068 48006
rect 15016 47942 15068 47948
rect 15028 47734 15056 47942
rect 15016 47728 15068 47734
rect 15016 47670 15068 47676
rect 15212 47036 15240 49166
rect 16040 49162 16068 52362
rect 16592 51406 16620 52498
rect 16776 52494 16804 53110
rect 16868 53106 16896 53926
rect 16960 53786 16988 53926
rect 16948 53780 17000 53786
rect 16948 53722 17000 53728
rect 17328 53446 17356 55694
rect 17684 55276 17736 55282
rect 17684 55218 17736 55224
rect 17696 54874 17724 55218
rect 17684 54868 17736 54874
rect 17684 54810 17736 54816
rect 17500 54528 17552 54534
rect 17500 54470 17552 54476
rect 17512 54126 17540 54470
rect 17500 54120 17552 54126
rect 17500 54062 17552 54068
rect 17972 54058 18000 57190
rect 18156 56846 18184 57326
rect 18248 56846 18276 61134
rect 19352 60858 19380 61746
rect 19616 61328 19668 61334
rect 19616 61270 19668 61276
rect 19432 61260 19484 61266
rect 19432 61202 19484 61208
rect 19340 60852 19392 60858
rect 19340 60794 19392 60800
rect 18788 60512 18840 60518
rect 18788 60454 18840 60460
rect 18800 60178 18828 60454
rect 19248 60240 19300 60246
rect 19248 60182 19300 60188
rect 18788 60172 18840 60178
rect 18788 60114 18840 60120
rect 18788 59628 18840 59634
rect 18788 59570 18840 59576
rect 18800 59430 18828 59570
rect 19260 59498 19288 60182
rect 19444 59770 19472 61202
rect 19628 61198 19656 61270
rect 19616 61192 19668 61198
rect 19616 61134 19668 61140
rect 19984 61056 20036 61062
rect 19984 60998 20036 61004
rect 19574 60956 19882 60976
rect 19574 60954 19580 60956
rect 19636 60954 19660 60956
rect 19716 60954 19740 60956
rect 19796 60954 19820 60956
rect 19876 60954 19882 60956
rect 19636 60902 19638 60954
rect 19818 60902 19820 60954
rect 19574 60900 19580 60902
rect 19636 60900 19660 60902
rect 19716 60900 19740 60902
rect 19796 60900 19820 60902
rect 19876 60900 19882 60902
rect 19574 60880 19882 60900
rect 19996 60722 20024 60998
rect 19984 60716 20036 60722
rect 19984 60658 20036 60664
rect 19984 60308 20036 60314
rect 19984 60250 20036 60256
rect 19574 59868 19882 59888
rect 19574 59866 19580 59868
rect 19636 59866 19660 59868
rect 19716 59866 19740 59868
rect 19796 59866 19820 59868
rect 19876 59866 19882 59868
rect 19636 59814 19638 59866
rect 19818 59814 19820 59866
rect 19574 59812 19580 59814
rect 19636 59812 19660 59814
rect 19716 59812 19740 59814
rect 19796 59812 19820 59814
rect 19876 59812 19882 59814
rect 19574 59792 19882 59812
rect 19432 59764 19484 59770
rect 19432 59706 19484 59712
rect 19524 59628 19576 59634
rect 19524 59570 19576 59576
rect 19248 59492 19300 59498
rect 19248 59434 19300 59440
rect 18788 59424 18840 59430
rect 18788 59366 18840 59372
rect 19064 58880 19116 58886
rect 19064 58822 19116 58828
rect 19076 58546 19104 58822
rect 19064 58540 19116 58546
rect 19064 58482 19116 58488
rect 19156 57792 19208 57798
rect 19156 57734 19208 57740
rect 19168 57458 19196 57734
rect 19156 57452 19208 57458
rect 19156 57394 19208 57400
rect 19260 57254 19288 59434
rect 19536 59158 19564 59570
rect 19996 59566 20024 60250
rect 19984 59560 20036 59566
rect 19984 59502 20036 59508
rect 19524 59152 19576 59158
rect 19524 59094 19576 59100
rect 19432 59016 19484 59022
rect 19432 58958 19484 58964
rect 19996 58970 20024 59502
rect 20168 59016 20220 59022
rect 19444 57934 19472 58958
rect 19996 58942 20116 58970
rect 20168 58958 20220 58964
rect 19984 58880 20036 58886
rect 19984 58822 20036 58828
rect 19574 58780 19882 58800
rect 19574 58778 19580 58780
rect 19636 58778 19660 58780
rect 19716 58778 19740 58780
rect 19796 58778 19820 58780
rect 19876 58778 19882 58780
rect 19636 58726 19638 58778
rect 19818 58726 19820 58778
rect 19574 58724 19580 58726
rect 19636 58724 19660 58726
rect 19716 58724 19740 58726
rect 19796 58724 19820 58726
rect 19876 58724 19882 58726
rect 19574 58704 19882 58724
rect 19996 58614 20024 58822
rect 19984 58608 20036 58614
rect 19984 58550 20036 58556
rect 19432 57928 19484 57934
rect 19432 57870 19484 57876
rect 19340 57588 19392 57594
rect 19340 57530 19392 57536
rect 19248 57248 19300 57254
rect 19248 57190 19300 57196
rect 18144 56840 18196 56846
rect 18144 56782 18196 56788
rect 18236 56840 18288 56846
rect 18236 56782 18288 56788
rect 18156 56234 18184 56782
rect 18144 56228 18196 56234
rect 18144 56170 18196 56176
rect 18248 55298 18276 56782
rect 19352 56166 19380 57530
rect 19444 56846 19472 57870
rect 19984 57792 20036 57798
rect 19984 57734 20036 57740
rect 19574 57692 19882 57712
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57616 19882 57636
rect 19996 57202 20024 57734
rect 20088 57390 20116 58942
rect 20180 58138 20208 58958
rect 20168 58132 20220 58138
rect 20168 58074 20220 58080
rect 20076 57384 20128 57390
rect 20076 57326 20128 57332
rect 19996 57174 20116 57202
rect 19432 56840 19484 56846
rect 19432 56782 19484 56788
rect 19984 56840 20036 56846
rect 19984 56782 20036 56788
rect 19432 56704 19484 56710
rect 19432 56646 19484 56652
rect 19444 56370 19472 56646
rect 19574 56604 19882 56624
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56528 19882 56548
rect 19432 56364 19484 56370
rect 19432 56306 19484 56312
rect 19340 56160 19392 56166
rect 19340 56102 19392 56108
rect 19352 55690 19380 56102
rect 19340 55684 19392 55690
rect 19340 55626 19392 55632
rect 19574 55516 19882 55536
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55440 19882 55460
rect 18156 55282 18276 55298
rect 18156 55276 18288 55282
rect 18156 55270 18236 55276
rect 18052 55072 18104 55078
rect 18052 55014 18104 55020
rect 18064 54126 18092 55014
rect 18052 54120 18104 54126
rect 18052 54062 18104 54068
rect 17960 54052 18012 54058
rect 17960 53994 18012 54000
rect 17408 53576 17460 53582
rect 17408 53518 17460 53524
rect 17316 53440 17368 53446
rect 17316 53382 17368 53388
rect 16856 53100 16908 53106
rect 16856 53042 16908 53048
rect 16764 52488 16816 52494
rect 16764 52430 16816 52436
rect 17132 52488 17184 52494
rect 17132 52430 17184 52436
rect 16580 51400 16632 51406
rect 16580 51342 16632 51348
rect 16764 51400 16816 51406
rect 16764 51342 16816 51348
rect 16776 51066 16804 51342
rect 16764 51060 16816 51066
rect 16764 51002 16816 51008
rect 16856 50924 16908 50930
rect 16856 50866 16908 50872
rect 16580 50176 16632 50182
rect 16580 50118 16632 50124
rect 16592 49162 16620 50118
rect 16868 49842 16896 50866
rect 16856 49836 16908 49842
rect 16856 49778 16908 49784
rect 16868 49722 16896 49778
rect 16776 49694 16896 49722
rect 16028 49156 16080 49162
rect 16028 49098 16080 49104
rect 16580 49156 16632 49162
rect 16580 49098 16632 49104
rect 16776 48142 16804 49694
rect 16856 49632 16908 49638
rect 16856 49574 16908 49580
rect 16868 49230 16896 49574
rect 16856 49224 16908 49230
rect 16856 49166 16908 49172
rect 17144 48754 17172 52430
rect 17328 50930 17356 53382
rect 17420 53242 17448 53518
rect 17408 53236 17460 53242
rect 17408 53178 17460 53184
rect 17592 52556 17644 52562
rect 17592 52498 17644 52504
rect 17408 51332 17460 51338
rect 17408 51274 17460 51280
rect 17420 51066 17448 51274
rect 17408 51060 17460 51066
rect 17408 51002 17460 51008
rect 17604 50930 17632 52498
rect 17972 52034 18000 53994
rect 18156 52494 18184 55270
rect 18236 55218 18288 55224
rect 19156 55072 19208 55078
rect 19156 55014 19208 55020
rect 19168 54670 19196 55014
rect 19996 54670 20024 56782
rect 20088 55622 20116 57174
rect 20076 55616 20128 55622
rect 20076 55558 20128 55564
rect 19156 54664 19208 54670
rect 19156 54606 19208 54612
rect 19984 54664 20036 54670
rect 19984 54606 20036 54612
rect 18236 54596 18288 54602
rect 18236 54538 18288 54544
rect 19248 54596 19300 54602
rect 19248 54538 19300 54544
rect 18248 54194 18276 54538
rect 19260 54262 19288 54538
rect 19340 54528 19392 54534
rect 19340 54470 19392 54476
rect 19432 54528 19484 54534
rect 19432 54470 19484 54476
rect 19248 54256 19300 54262
rect 19248 54198 19300 54204
rect 18236 54188 18288 54194
rect 18236 54130 18288 54136
rect 18328 54120 18380 54126
rect 18328 54062 18380 54068
rect 18512 54120 18564 54126
rect 18564 54080 18644 54108
rect 18512 54062 18564 54068
rect 18340 53990 18368 54062
rect 18328 53984 18380 53990
rect 18328 53926 18380 53932
rect 18616 53446 18644 54080
rect 19352 53990 19380 54470
rect 19444 54194 19472 54470
rect 19574 54428 19882 54448
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54352 19882 54372
rect 19432 54188 19484 54194
rect 19432 54130 19484 54136
rect 19340 53984 19392 53990
rect 19340 53926 19392 53932
rect 19352 53514 19380 53926
rect 18880 53508 18932 53514
rect 18880 53450 18932 53456
rect 19340 53508 19392 53514
rect 19340 53450 19392 53456
rect 18604 53440 18656 53446
rect 18604 53382 18656 53388
rect 18052 52488 18104 52494
rect 18052 52430 18104 52436
rect 18144 52488 18196 52494
rect 18144 52430 18196 52436
rect 17880 52006 18000 52034
rect 17880 51814 17908 52006
rect 18064 51898 18092 52430
rect 17972 51882 18092 51898
rect 17960 51876 18092 51882
rect 18012 51870 18092 51876
rect 17960 51818 18012 51824
rect 17868 51808 17920 51814
rect 17920 51756 18000 51762
rect 17868 51750 18000 51756
rect 17880 51734 18000 51750
rect 17972 51542 18000 51734
rect 18064 51610 18092 51870
rect 18052 51604 18104 51610
rect 18052 51546 18104 51552
rect 17960 51536 18012 51542
rect 17960 51478 18012 51484
rect 18156 51474 18184 52430
rect 18328 52420 18380 52426
rect 18328 52362 18380 52368
rect 18340 52018 18368 52362
rect 18328 52012 18380 52018
rect 18328 51954 18380 51960
rect 18616 51950 18644 53382
rect 18420 51944 18472 51950
rect 18420 51886 18472 51892
rect 18604 51944 18656 51950
rect 18604 51886 18656 51892
rect 18144 51468 18196 51474
rect 18144 51410 18196 51416
rect 18432 51406 18460 51886
rect 18420 51400 18472 51406
rect 18420 51342 18472 51348
rect 17316 50924 17368 50930
rect 17316 50866 17368 50872
rect 17592 50924 17644 50930
rect 17592 50866 17644 50872
rect 18512 50312 18564 50318
rect 18512 50254 18564 50260
rect 17684 50176 17736 50182
rect 17684 50118 17736 50124
rect 17696 49978 17724 50118
rect 17684 49972 17736 49978
rect 17684 49914 17736 49920
rect 17592 49768 17644 49774
rect 17592 49710 17644 49716
rect 17604 49434 17632 49710
rect 18236 49700 18288 49706
rect 18236 49642 18288 49648
rect 17592 49428 17644 49434
rect 17592 49370 17644 49376
rect 17316 49224 17368 49230
rect 17316 49166 17368 49172
rect 17132 48748 17184 48754
rect 17132 48690 17184 48696
rect 15292 48136 15344 48142
rect 15292 48078 15344 48084
rect 16764 48136 16816 48142
rect 16764 48078 16816 48084
rect 15304 47258 15332 48078
rect 16304 48000 16356 48006
rect 16304 47942 16356 47948
rect 17040 48000 17092 48006
rect 17040 47942 17092 47948
rect 15568 47524 15620 47530
rect 15568 47466 15620 47472
rect 15292 47252 15344 47258
rect 15292 47194 15344 47200
rect 15580 47122 15608 47466
rect 16316 47122 16344 47942
rect 15568 47116 15620 47122
rect 15568 47058 15620 47064
rect 16304 47116 16356 47122
rect 16304 47058 16356 47064
rect 17052 47054 17080 47942
rect 17328 47666 17356 49166
rect 17408 48136 17460 48142
rect 17408 48078 17460 48084
rect 17420 47802 17448 48078
rect 17960 48068 18012 48074
rect 17960 48010 18012 48016
rect 18052 48068 18104 48074
rect 18052 48010 18104 48016
rect 17972 47802 18000 48010
rect 17408 47796 17460 47802
rect 17408 47738 17460 47744
rect 17960 47796 18012 47802
rect 17960 47738 18012 47744
rect 18064 47666 18092 48010
rect 17316 47660 17368 47666
rect 17316 47602 17368 47608
rect 18052 47660 18104 47666
rect 18052 47602 18104 47608
rect 15292 47048 15344 47054
rect 15212 47008 15292 47036
rect 15292 46990 15344 46996
rect 17040 47048 17092 47054
rect 17040 46990 17092 46996
rect 15200 45824 15252 45830
rect 15200 45766 15252 45772
rect 15212 45558 15240 45766
rect 15200 45552 15252 45558
rect 15200 45494 15252 45500
rect 15304 44878 15332 46990
rect 17328 46646 17356 47602
rect 17684 47592 17736 47598
rect 17684 47534 17736 47540
rect 17696 47258 17724 47534
rect 18248 47530 18276 49642
rect 18524 49434 18552 50254
rect 18604 50244 18656 50250
rect 18604 50186 18656 50192
rect 18616 49842 18644 50186
rect 18604 49836 18656 49842
rect 18604 49778 18656 49784
rect 18892 49586 18920 53450
rect 19574 53340 19882 53360
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53264 19882 53284
rect 19996 53106 20024 54606
rect 20088 53514 20116 55558
rect 20168 54528 20220 54534
rect 20168 54470 20220 54476
rect 20180 54262 20208 54470
rect 20168 54256 20220 54262
rect 20168 54198 20220 54204
rect 20076 53508 20128 53514
rect 20076 53450 20128 53456
rect 20168 53508 20220 53514
rect 20168 53450 20220 53456
rect 19984 53100 20036 53106
rect 19984 53042 20036 53048
rect 19340 52896 19392 52902
rect 19340 52838 19392 52844
rect 19352 52562 19380 52838
rect 19340 52556 19392 52562
rect 19340 52498 19392 52504
rect 19432 52420 19484 52426
rect 19432 52362 19484 52368
rect 18972 51944 19024 51950
rect 18972 51886 19024 51892
rect 18984 49774 19012 51886
rect 19248 51808 19300 51814
rect 19248 51750 19300 51756
rect 19260 51542 19288 51750
rect 19444 51610 19472 52362
rect 19574 52252 19882 52272
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52176 19882 52196
rect 20088 52086 20116 53450
rect 20076 52080 20128 52086
rect 20076 52022 20128 52028
rect 20180 51950 20208 53450
rect 20168 51944 20220 51950
rect 20168 51886 20220 51892
rect 19892 51808 19944 51814
rect 20076 51808 20128 51814
rect 19944 51768 20024 51796
rect 19892 51750 19944 51756
rect 19432 51604 19484 51610
rect 19432 51546 19484 51552
rect 19248 51536 19300 51542
rect 19248 51478 19300 51484
rect 19574 51164 19882 51184
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51088 19882 51108
rect 19996 51074 20024 51768
rect 20076 51750 20128 51756
rect 20088 51406 20116 51750
rect 20076 51400 20128 51406
rect 20076 51342 20128 51348
rect 20272 51074 20300 69226
rect 20720 61804 20772 61810
rect 20720 61746 20772 61752
rect 20352 61600 20404 61606
rect 20352 61542 20404 61548
rect 20364 61402 20392 61542
rect 20732 61402 20760 61746
rect 21088 61600 21140 61606
rect 21088 61542 21140 61548
rect 21180 61600 21232 61606
rect 21180 61542 21232 61548
rect 20352 61396 20404 61402
rect 20352 61338 20404 61344
rect 20720 61396 20772 61402
rect 20720 61338 20772 61344
rect 21100 61198 21128 61542
rect 21192 61266 21220 61542
rect 21180 61260 21232 61266
rect 21180 61202 21232 61208
rect 21088 61192 21140 61198
rect 21088 61134 21140 61140
rect 20812 61056 20864 61062
rect 20812 60998 20864 61004
rect 20824 60178 20852 60998
rect 21548 60512 21600 60518
rect 21548 60454 21600 60460
rect 21560 60178 21588 60454
rect 20812 60172 20864 60178
rect 20812 60114 20864 60120
rect 21548 60172 21600 60178
rect 21548 60114 21600 60120
rect 20996 60104 21048 60110
rect 20996 60046 21048 60052
rect 20352 59424 20404 59430
rect 20352 59366 20404 59372
rect 20364 58682 20392 59366
rect 20444 58948 20496 58954
rect 20444 58890 20496 58896
rect 20352 58676 20404 58682
rect 20352 58618 20404 58624
rect 20364 57866 20392 58618
rect 20456 58342 20484 58890
rect 20628 58676 20680 58682
rect 20628 58618 20680 58624
rect 20444 58336 20496 58342
rect 20444 58278 20496 58284
rect 20456 58070 20484 58278
rect 20444 58064 20496 58070
rect 20444 58006 20496 58012
rect 20352 57860 20404 57866
rect 20352 57802 20404 57808
rect 20352 56704 20404 56710
rect 20352 56646 20404 56652
rect 20364 56438 20392 56646
rect 20352 56432 20404 56438
rect 20352 56374 20404 56380
rect 20456 55894 20484 58006
rect 20640 57798 20668 58618
rect 21008 58614 21036 60046
rect 21272 59016 21324 59022
rect 21272 58958 21324 58964
rect 21284 58682 21312 58958
rect 21456 58880 21508 58886
rect 21456 58822 21508 58828
rect 21272 58676 21324 58682
rect 21272 58618 21324 58624
rect 21468 58614 21496 58822
rect 20996 58608 21048 58614
rect 20996 58550 21048 58556
rect 21456 58608 21508 58614
rect 21456 58550 21508 58556
rect 20996 58472 21048 58478
rect 20996 58414 21048 58420
rect 21008 58138 21036 58414
rect 20996 58132 21048 58138
rect 20996 58074 21048 58080
rect 20628 57792 20680 57798
rect 20628 57734 20680 57740
rect 20536 56840 20588 56846
rect 20536 56782 20588 56788
rect 20548 55962 20576 56782
rect 20536 55956 20588 55962
rect 20536 55898 20588 55904
rect 20444 55888 20496 55894
rect 20444 55830 20496 55836
rect 20352 54664 20404 54670
rect 20352 54606 20404 54612
rect 20364 53786 20392 54606
rect 20352 53780 20404 53786
rect 20352 53722 20404 53728
rect 20456 53718 20484 55830
rect 20628 54120 20680 54126
rect 20628 54062 20680 54068
rect 20444 53712 20496 53718
rect 20444 53654 20496 53660
rect 20352 52080 20404 52086
rect 20352 52022 20404 52028
rect 20364 51406 20392 52022
rect 20352 51400 20404 51406
rect 20352 51342 20404 51348
rect 19996 51046 20116 51074
rect 20272 51046 20392 51074
rect 20456 51066 20484 53654
rect 20536 51332 20588 51338
rect 20536 51274 20588 51280
rect 19524 50720 19576 50726
rect 19524 50662 19576 50668
rect 19536 50318 19564 50662
rect 20088 50318 20116 51046
rect 20260 50924 20312 50930
rect 20260 50866 20312 50872
rect 19340 50312 19392 50318
rect 19340 50254 19392 50260
rect 19524 50312 19576 50318
rect 19524 50254 19576 50260
rect 20076 50312 20128 50318
rect 20076 50254 20128 50260
rect 18972 49768 19024 49774
rect 19024 49716 19104 49722
rect 18972 49710 19104 49716
rect 18984 49694 19104 49710
rect 18892 49558 19012 49586
rect 18512 49428 18564 49434
rect 18512 49370 18564 49376
rect 18880 47592 18932 47598
rect 18880 47534 18932 47540
rect 18236 47524 18288 47530
rect 18236 47466 18288 47472
rect 17684 47252 17736 47258
rect 17684 47194 17736 47200
rect 17316 46640 17368 46646
rect 17316 46582 17368 46588
rect 17408 46572 17460 46578
rect 17408 46514 17460 46520
rect 17500 46572 17552 46578
rect 17500 46514 17552 46520
rect 17420 46170 17448 46514
rect 17408 46164 17460 46170
rect 17408 46106 17460 46112
rect 15476 45960 15528 45966
rect 15476 45902 15528 45908
rect 16580 45960 16632 45966
rect 16580 45902 16632 45908
rect 15488 45082 15516 45902
rect 16592 45626 16620 45902
rect 16580 45620 16632 45626
rect 16580 45562 16632 45568
rect 17420 45490 17448 46106
rect 16948 45484 17000 45490
rect 16948 45426 17000 45432
rect 17408 45484 17460 45490
rect 17408 45426 17460 45432
rect 15936 45280 15988 45286
rect 15936 45222 15988 45228
rect 15476 45076 15528 45082
rect 15476 45018 15528 45024
rect 15948 44946 15976 45222
rect 15936 44940 15988 44946
rect 15936 44882 15988 44888
rect 15292 44872 15344 44878
rect 15292 44814 15344 44820
rect 15568 44872 15620 44878
rect 15568 44814 15620 44820
rect 15384 44396 15436 44402
rect 15384 44338 15436 44344
rect 15200 44192 15252 44198
rect 15200 44134 15252 44140
rect 15212 43790 15240 44134
rect 15200 43784 15252 43790
rect 15200 43726 15252 43732
rect 15396 43450 15424 44338
rect 15384 43444 15436 43450
rect 15384 43386 15436 43392
rect 15580 43314 15608 44814
rect 16764 44260 16816 44266
rect 16764 44202 16816 44208
rect 16776 43926 16804 44202
rect 16856 44192 16908 44198
rect 16856 44134 16908 44140
rect 16580 43920 16632 43926
rect 16580 43862 16632 43868
rect 16764 43920 16816 43926
rect 16764 43862 16816 43868
rect 15752 43716 15804 43722
rect 15752 43658 15804 43664
rect 15764 43450 15792 43658
rect 15752 43444 15804 43450
rect 15752 43386 15804 43392
rect 16592 43382 16620 43862
rect 16868 43790 16896 44134
rect 16856 43784 16908 43790
rect 16856 43726 16908 43732
rect 16764 43648 16816 43654
rect 16764 43590 16816 43596
rect 16580 43376 16632 43382
rect 16580 43318 16632 43324
rect 16776 43314 16804 43590
rect 15568 43308 15620 43314
rect 15568 43250 15620 43256
rect 16764 43308 16816 43314
rect 16764 43250 16816 43256
rect 15476 42560 15528 42566
rect 15476 42502 15528 42508
rect 15488 42294 15516 42502
rect 15476 42288 15528 42294
rect 15476 42230 15528 42236
rect 14832 41744 14884 41750
rect 14832 41686 14884 41692
rect 15580 41614 15608 43250
rect 16960 42702 16988 45426
rect 17040 44396 17092 44402
rect 17040 44338 17092 44344
rect 17052 43450 17080 44338
rect 17040 43444 17092 43450
rect 17040 43386 17092 43392
rect 17512 42702 17540 46514
rect 18248 45354 18276 47466
rect 18892 47462 18920 47534
rect 18880 47456 18932 47462
rect 18880 47398 18932 47404
rect 18984 46578 19012 49558
rect 19076 47598 19104 49694
rect 19352 49434 19380 50254
rect 19984 50176 20036 50182
rect 19984 50118 20036 50124
rect 19574 50076 19882 50096
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50000 19882 50020
rect 19996 49978 20024 50118
rect 19984 49972 20036 49978
rect 19984 49914 20036 49920
rect 20088 49638 20116 50254
rect 20272 49978 20300 50866
rect 20260 49972 20312 49978
rect 20260 49914 20312 49920
rect 20260 49836 20312 49842
rect 20260 49778 20312 49784
rect 20076 49632 20128 49638
rect 20076 49574 20128 49580
rect 19340 49428 19392 49434
rect 19340 49370 19392 49376
rect 19574 48988 19882 49008
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48912 19882 48932
rect 20088 48872 20116 49574
rect 20272 49314 20300 49778
rect 19812 48844 20116 48872
rect 19812 48346 19840 48844
rect 19984 48748 20036 48754
rect 19984 48690 20036 48696
rect 19996 48346 20024 48690
rect 19800 48340 19852 48346
rect 19800 48282 19852 48288
rect 19984 48340 20036 48346
rect 19984 48282 20036 48288
rect 19574 47900 19882 47920
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47824 19882 47844
rect 19064 47592 19116 47598
rect 19064 47534 19116 47540
rect 18972 46572 19024 46578
rect 18972 46514 19024 46520
rect 18512 46368 18564 46374
rect 18512 46310 18564 46316
rect 18524 45966 18552 46310
rect 18984 45966 19012 46514
rect 18512 45960 18564 45966
rect 18512 45902 18564 45908
rect 18972 45960 19024 45966
rect 18972 45902 19024 45908
rect 18420 45484 18472 45490
rect 18420 45426 18472 45432
rect 18236 45348 18288 45354
rect 18236 45290 18288 45296
rect 18248 44418 18276 45290
rect 18432 45286 18460 45426
rect 19076 45422 19104 47534
rect 19984 46912 20036 46918
rect 19984 46854 20036 46860
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19996 46578 20024 46854
rect 19984 46572 20036 46578
rect 19984 46514 20036 46520
rect 19248 46368 19300 46374
rect 19248 46310 19300 46316
rect 19708 46368 19760 46374
rect 19708 46310 19760 46316
rect 19260 46050 19288 46310
rect 19168 46034 19288 46050
rect 19168 46028 19300 46034
rect 19168 46022 19248 46028
rect 19064 45416 19116 45422
rect 19064 45358 19116 45364
rect 18420 45280 18472 45286
rect 18420 45222 18472 45228
rect 18248 44390 18368 44418
rect 17960 44328 18012 44334
rect 17960 44270 18012 44276
rect 17972 42770 18000 44270
rect 18340 44266 18368 44390
rect 19168 44334 19196 46022
rect 19248 45970 19300 45976
rect 19720 45898 19748 46310
rect 19984 46164 20036 46170
rect 20088 46152 20116 48844
rect 20180 49286 20300 49314
rect 20180 48006 20208 49286
rect 20260 49156 20312 49162
rect 20260 49098 20312 49104
rect 20272 48754 20300 49098
rect 20260 48748 20312 48754
rect 20260 48690 20312 48696
rect 20168 48000 20220 48006
rect 20168 47942 20220 47948
rect 20180 47122 20208 47942
rect 20168 47116 20220 47122
rect 20168 47058 20220 47064
rect 20036 46124 20116 46152
rect 19984 46106 20036 46112
rect 20180 45898 20208 47058
rect 19248 45892 19300 45898
rect 19248 45834 19300 45840
rect 19708 45892 19760 45898
rect 19708 45834 19760 45840
rect 20168 45892 20220 45898
rect 20168 45834 20220 45840
rect 19260 45626 19288 45834
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19248 45620 19300 45626
rect 19248 45562 19300 45568
rect 20076 45484 20128 45490
rect 20076 45426 20128 45432
rect 19432 45416 19484 45422
rect 19432 45358 19484 45364
rect 19444 45082 19472 45358
rect 20088 45082 20116 45426
rect 19432 45076 19484 45082
rect 19432 45018 19484 45024
rect 20076 45076 20128 45082
rect 20076 45018 20128 45024
rect 19892 45008 19944 45014
rect 19944 44956 20116 44962
rect 19892 44950 20116 44956
rect 19904 44934 20116 44950
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 18972 44328 19024 44334
rect 18972 44270 19024 44276
rect 19156 44328 19208 44334
rect 19156 44270 19208 44276
rect 18328 44260 18380 44266
rect 18328 44202 18380 44208
rect 18340 43926 18368 44202
rect 18328 43920 18380 43926
rect 18328 43862 18380 43868
rect 18984 43178 19012 44270
rect 19064 43920 19116 43926
rect 19064 43862 19116 43868
rect 19076 43178 19104 43862
rect 19168 43450 19196 44270
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19156 43444 19208 43450
rect 19156 43386 19208 43392
rect 19340 43240 19392 43246
rect 19340 43182 19392 43188
rect 18972 43172 19024 43178
rect 18972 43114 19024 43120
rect 19064 43172 19116 43178
rect 19064 43114 19116 43120
rect 17960 42764 18012 42770
rect 17960 42706 18012 42712
rect 15752 42696 15804 42702
rect 15752 42638 15804 42644
rect 16948 42696 17000 42702
rect 16948 42638 17000 42644
rect 17500 42696 17552 42702
rect 17500 42638 17552 42644
rect 17972 42650 18000 42706
rect 15764 41818 15792 42638
rect 16948 42560 17000 42566
rect 16948 42502 17000 42508
rect 16960 42226 16988 42502
rect 17512 42294 17540 42638
rect 17972 42622 18092 42650
rect 17960 42560 18012 42566
rect 17960 42502 18012 42508
rect 17500 42288 17552 42294
rect 17500 42230 17552 42236
rect 16948 42220 17000 42226
rect 16948 42162 17000 42168
rect 17224 42220 17276 42226
rect 17224 42162 17276 42168
rect 16120 42016 16172 42022
rect 16120 41958 16172 41964
rect 15752 41812 15804 41818
rect 15752 41754 15804 41760
rect 16132 41682 16160 41958
rect 16120 41676 16172 41682
rect 16120 41618 16172 41624
rect 15568 41608 15620 41614
rect 15568 41550 15620 41556
rect 17236 41274 17264 42162
rect 17592 41608 17644 41614
rect 17592 41550 17644 41556
rect 17224 41268 17276 41274
rect 17224 41210 17276 41216
rect 14464 35760 14516 35766
rect 14464 35702 14516 35708
rect 8024 35556 8076 35562
rect 8024 35498 8076 35504
rect 14476 35494 14504 35702
rect 14464 35488 14516 35494
rect 14464 35430 14516 35436
rect 13820 27940 13872 27946
rect 13820 27882 13872 27888
rect 13832 16574 13860 27882
rect 13832 16546 14872 16574
rect 10232 4548 10284 4554
rect 10232 4490 10284 4496
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4632 3602 4660 3878
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4618 3496 4674 3505
rect 5184 3466 5212 3878
rect 4618 3431 4674 3440
rect 5172 3460 5224 3466
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3252 800 3280 2382
rect 4632 1714 4660 3431
rect 5172 3402 5224 3408
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 4540 1686 4660 1714
rect 4540 800 4568 1686
rect 5828 800 5856 2518
rect 6564 2514 6592 3334
rect 6656 3058 6684 3402
rect 6840 3126 6868 3878
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 10244 3058 10272 4490
rect 13542 3632 13598 3641
rect 10968 3596 11020 3602
rect 13542 3567 13598 3576
rect 10968 3538 11020 3544
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 7116 800 7144 2926
rect 10428 2650 10456 3470
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10612 3126 10640 3402
rect 10600 3120 10652 3126
rect 10600 3062 10652 3068
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10980 800 11008 3538
rect 13556 800 13584 3567
rect 14844 800 14872 16546
rect 17604 7750 17632 41550
rect 17684 41540 17736 41546
rect 17684 41482 17736 41488
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17696 2650 17724 41482
rect 17972 41138 18000 42502
rect 18064 42362 18092 42622
rect 18788 42628 18840 42634
rect 18788 42570 18840 42576
rect 18052 42356 18104 42362
rect 18052 42298 18104 42304
rect 18420 42356 18472 42362
rect 18420 42298 18472 42304
rect 18432 41750 18460 42298
rect 18800 42226 18828 42570
rect 19352 42226 19380 43182
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 18788 42220 18840 42226
rect 18788 42162 18840 42168
rect 19340 42220 19392 42226
rect 19340 42162 19392 42168
rect 19616 42220 19668 42226
rect 19616 42162 19668 42168
rect 19248 42016 19300 42022
rect 19248 41958 19300 41964
rect 18420 41744 18472 41750
rect 18420 41686 18472 41692
rect 19260 41682 19288 41958
rect 19628 41818 19656 42162
rect 19984 42016 20036 42022
rect 19984 41958 20036 41964
rect 19616 41812 19668 41818
rect 19616 41754 19668 41760
rect 19248 41676 19300 41682
rect 19248 41618 19300 41624
rect 19432 41472 19484 41478
rect 19432 41414 19484 41420
rect 19444 41274 19472 41414
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19432 41268 19484 41274
rect 19432 41210 19484 41216
rect 19996 41138 20024 41958
rect 17960 41132 18012 41138
rect 17960 41074 18012 41080
rect 19984 41132 20036 41138
rect 19984 41074 20036 41080
rect 19248 41064 19300 41070
rect 19248 41006 19300 41012
rect 19260 40594 19288 41006
rect 19248 40588 19300 40594
rect 19248 40530 19300 40536
rect 19984 40384 20036 40390
rect 19984 40326 20036 40332
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19996 40050 20024 40326
rect 19984 40044 20036 40050
rect 19984 39986 20036 39992
rect 19432 39296 19484 39302
rect 19432 39238 19484 39244
rect 19444 39098 19472 39238
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19432 39092 19484 39098
rect 19432 39034 19484 39040
rect 19996 38962 20024 39986
rect 19984 38956 20036 38962
rect 19984 38898 20036 38904
rect 19996 38350 20024 38898
rect 19984 38344 20036 38350
rect 19984 38286 20036 38292
rect 19984 38208 20036 38214
rect 19984 38150 20036 38156
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19996 37942 20024 38150
rect 19984 37936 20036 37942
rect 19984 37878 20036 37884
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19156 35692 19208 35698
rect 19156 35634 19208 35640
rect 19984 35692 20036 35698
rect 19984 35634 20036 35640
rect 19168 21350 19196 35634
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19156 21344 19208 21350
rect 19156 21286 19208 21292
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19996 7818 20024 35634
rect 20088 35290 20116 44934
rect 20260 43648 20312 43654
rect 20260 43590 20312 43596
rect 20272 43314 20300 43590
rect 20260 43308 20312 43314
rect 20260 43250 20312 43256
rect 20168 43240 20220 43246
rect 20168 43182 20220 43188
rect 20180 42090 20208 43182
rect 20168 42084 20220 42090
rect 20168 42026 20220 42032
rect 20364 35630 20392 51046
rect 20444 51060 20496 51066
rect 20444 51002 20496 51008
rect 20548 49230 20576 51274
rect 20640 49774 20668 54062
rect 20904 53100 20956 53106
rect 20904 53042 20956 53048
rect 20720 52352 20772 52358
rect 20720 52294 20772 52300
rect 20732 52018 20760 52294
rect 20720 52012 20772 52018
rect 20720 51954 20772 51960
rect 20628 49768 20680 49774
rect 20628 49710 20680 49716
rect 20536 49224 20588 49230
rect 20536 49166 20588 49172
rect 20548 48686 20576 49166
rect 20720 48884 20772 48890
rect 20720 48826 20772 48832
rect 20536 48680 20588 48686
rect 20536 48622 20588 48628
rect 20444 48544 20496 48550
rect 20444 48486 20496 48492
rect 20456 48210 20484 48486
rect 20444 48204 20496 48210
rect 20444 48146 20496 48152
rect 20732 48142 20760 48826
rect 20812 48816 20864 48822
rect 20812 48758 20864 48764
rect 20720 48136 20772 48142
rect 20720 48078 20772 48084
rect 20824 47054 20852 48758
rect 20916 48736 20944 53042
rect 21364 52420 21416 52426
rect 21364 52362 21416 52368
rect 21376 52086 21404 52362
rect 21364 52080 21416 52086
rect 21364 52022 21416 52028
rect 20996 50924 21048 50930
rect 20996 50866 21048 50872
rect 21008 50454 21036 50866
rect 20996 50448 21048 50454
rect 20996 50390 21048 50396
rect 21652 50402 21680 69226
rect 21824 62280 21876 62286
rect 21824 62222 21876 62228
rect 21836 61810 21864 62222
rect 21824 61804 21876 61810
rect 21824 61746 21876 61752
rect 22008 60648 22060 60654
rect 22008 60590 22060 60596
rect 21732 60104 21784 60110
rect 22020 60058 22048 60590
rect 21784 60052 22048 60058
rect 21732 60046 22048 60052
rect 21744 60030 22048 60046
rect 22020 59430 22048 60030
rect 22008 59424 22060 59430
rect 22008 59366 22060 59372
rect 21732 56840 21784 56846
rect 21732 56782 21784 56788
rect 21744 56370 21772 56782
rect 21732 56364 21784 56370
rect 21732 56306 21784 56312
rect 21744 54738 21772 56306
rect 21824 54800 21876 54806
rect 21824 54742 21876 54748
rect 21732 54732 21784 54738
rect 21732 54674 21784 54680
rect 21744 54194 21772 54674
rect 21732 54188 21784 54194
rect 21732 54130 21784 54136
rect 21744 53582 21772 54130
rect 21732 53576 21784 53582
rect 21732 53518 21784 53524
rect 21744 53106 21772 53518
rect 21732 53100 21784 53106
rect 21732 53042 21784 53048
rect 21732 52964 21784 52970
rect 21732 52906 21784 52912
rect 21744 52630 21772 52906
rect 21732 52624 21784 52630
rect 21732 52566 21784 52572
rect 21836 52494 21864 54742
rect 21916 54596 21968 54602
rect 21916 54538 21968 54544
rect 21928 54262 21956 54538
rect 21916 54256 21968 54262
rect 21916 54198 21968 54204
rect 21824 52488 21876 52494
rect 21824 52430 21876 52436
rect 21824 51536 21876 51542
rect 21824 51478 21876 51484
rect 21456 50380 21508 50386
rect 21652 50374 21772 50402
rect 21456 50322 21508 50328
rect 20996 48748 21048 48754
rect 20916 48708 20996 48736
rect 20996 48690 21048 48696
rect 21008 47598 21036 48690
rect 20996 47592 21048 47598
rect 20996 47534 21048 47540
rect 21088 47456 21140 47462
rect 21088 47398 21140 47404
rect 20812 47048 20864 47054
rect 20996 47048 21048 47054
rect 20864 46996 20944 47002
rect 20812 46990 20944 46996
rect 20996 46990 21048 46996
rect 20824 46974 20944 46990
rect 20812 46912 20864 46918
rect 20812 46854 20864 46860
rect 20824 46646 20852 46854
rect 20812 46640 20864 46646
rect 20812 46582 20864 46588
rect 20916 46578 20944 46974
rect 20904 46572 20956 46578
rect 20904 46514 20956 46520
rect 20916 46458 20944 46514
rect 20824 46430 20944 46458
rect 20536 45892 20588 45898
rect 20536 45834 20588 45840
rect 20548 45286 20576 45834
rect 20628 45824 20680 45830
rect 20628 45766 20680 45772
rect 20640 45626 20668 45766
rect 20628 45620 20680 45626
rect 20628 45562 20680 45568
rect 20536 45280 20588 45286
rect 20536 45222 20588 45228
rect 20548 44538 20576 45222
rect 20824 44946 20852 46430
rect 21008 46102 21036 46990
rect 20996 46096 21048 46102
rect 20996 46038 21048 46044
rect 20904 45824 20956 45830
rect 20904 45766 20956 45772
rect 20812 44940 20864 44946
rect 20812 44882 20864 44888
rect 20916 44878 20944 45766
rect 21100 44946 21128 47398
rect 21364 45552 21416 45558
rect 21364 45494 21416 45500
rect 21272 45484 21324 45490
rect 21272 45426 21324 45432
rect 21088 44940 21140 44946
rect 21088 44882 21140 44888
rect 20904 44872 20956 44878
rect 20904 44814 20956 44820
rect 20720 44804 20772 44810
rect 20720 44746 20772 44752
rect 20536 44532 20588 44538
rect 20536 44474 20588 44480
rect 20536 43988 20588 43994
rect 20536 43930 20588 43936
rect 20548 43450 20576 43930
rect 20732 43722 20760 44746
rect 20996 44192 21048 44198
rect 20996 44134 21048 44140
rect 21008 43858 21036 44134
rect 20996 43852 21048 43858
rect 20996 43794 21048 43800
rect 21180 43784 21232 43790
rect 21180 43726 21232 43732
rect 20720 43716 20772 43722
rect 20720 43658 20772 43664
rect 21088 43648 21140 43654
rect 21088 43590 21140 43596
rect 20444 43444 20496 43450
rect 20444 43386 20496 43392
rect 20536 43444 20588 43450
rect 20536 43386 20588 43392
rect 20456 43246 20484 43386
rect 20444 43240 20496 43246
rect 20444 43182 20496 43188
rect 20996 42628 21048 42634
rect 20996 42570 21048 42576
rect 21008 42226 21036 42570
rect 20996 42220 21048 42226
rect 20996 42162 21048 42168
rect 20720 39364 20772 39370
rect 20720 39306 20772 39312
rect 20732 38554 20760 39306
rect 21100 38962 21128 43590
rect 21192 43246 21220 43726
rect 21180 43240 21232 43246
rect 21180 43182 21232 43188
rect 21192 42770 21220 43182
rect 21284 43178 21312 45426
rect 21376 43790 21404 45494
rect 21468 45082 21496 50322
rect 21640 46368 21692 46374
rect 21640 46310 21692 46316
rect 21652 46034 21680 46310
rect 21640 46028 21692 46034
rect 21640 45970 21692 45976
rect 21640 45824 21692 45830
rect 21640 45766 21692 45772
rect 21652 45490 21680 45766
rect 21640 45484 21692 45490
rect 21640 45426 21692 45432
rect 21456 45076 21508 45082
rect 21456 45018 21508 45024
rect 21364 43784 21416 43790
rect 21364 43726 21416 43732
rect 21548 43648 21600 43654
rect 21548 43590 21600 43596
rect 21272 43172 21324 43178
rect 21272 43114 21324 43120
rect 21180 42764 21232 42770
rect 21180 42706 21232 42712
rect 21560 42566 21588 43590
rect 21640 43104 21692 43110
rect 21640 43046 21692 43052
rect 21652 42702 21680 43046
rect 21640 42696 21692 42702
rect 21640 42638 21692 42644
rect 21548 42560 21600 42566
rect 21548 42502 21600 42508
rect 21180 41608 21232 41614
rect 21178 41576 21180 41585
rect 21232 41576 21234 41585
rect 21178 41511 21234 41520
rect 21272 40520 21324 40526
rect 21272 40462 21324 40468
rect 21284 39846 21312 40462
rect 21548 40384 21600 40390
rect 21548 40326 21600 40332
rect 21560 40050 21588 40326
rect 21548 40044 21600 40050
rect 21548 39986 21600 39992
rect 21272 39840 21324 39846
rect 21272 39782 21324 39788
rect 21284 39506 21312 39782
rect 21272 39500 21324 39506
rect 21272 39442 21324 39448
rect 20904 38956 20956 38962
rect 20904 38898 20956 38904
rect 21088 38956 21140 38962
rect 21088 38898 21140 38904
rect 20720 38548 20772 38554
rect 20720 38490 20772 38496
rect 20916 38214 20944 38898
rect 21180 38752 21232 38758
rect 21180 38694 21232 38700
rect 21192 38282 21220 38694
rect 21180 38276 21232 38282
rect 21180 38218 21232 38224
rect 20904 38208 20956 38214
rect 20904 38150 20956 38156
rect 20916 38010 20944 38150
rect 20904 38004 20956 38010
rect 20904 37946 20956 37952
rect 20720 35692 20772 35698
rect 20720 35634 20772 35640
rect 20352 35624 20404 35630
rect 20352 35566 20404 35572
rect 20076 35284 20128 35290
rect 20076 35226 20128 35232
rect 20536 35012 20588 35018
rect 20536 34954 20588 34960
rect 20548 34610 20576 34954
rect 20536 34604 20588 34610
rect 20536 34546 20588 34552
rect 20732 24614 20760 35634
rect 20904 35624 20956 35630
rect 20904 35566 20956 35572
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20720 24608 20772 24614
rect 20720 24550 20772 24556
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19352 3058 19380 3470
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19524 2984 19576 2990
rect 19524 2926 19576 2932
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19536 2650 19564 2926
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17420 800 17448 2382
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2926
rect 20824 2310 20852 35022
rect 20916 2378 20944 35566
rect 21744 35290 21772 50374
rect 21836 47054 21864 51478
rect 21824 47048 21876 47054
rect 21824 46990 21876 46996
rect 22112 46714 22140 71318
rect 23174 71200 23286 71318
rect 23818 71200 23930 72000
rect 25106 71200 25218 72000
rect 26394 71200 26506 72000
rect 27682 71200 27794 72000
rect 28970 71346 29082 72000
rect 28970 71318 29408 71346
rect 28970 71200 29082 71318
rect 24860 69216 24912 69222
rect 24860 69158 24912 69164
rect 24872 68882 24900 69158
rect 25148 68882 25176 71200
rect 27344 69216 27396 69222
rect 27344 69158 27396 69164
rect 27356 68882 27384 69158
rect 27724 68882 27752 71200
rect 24860 68876 24912 68882
rect 24860 68818 24912 68824
rect 25136 68876 25188 68882
rect 25136 68818 25188 68824
rect 27344 68876 27396 68882
rect 27344 68818 27396 68824
rect 27712 68876 27764 68882
rect 27712 68818 27764 68824
rect 24860 68740 24912 68746
rect 24860 68682 24912 68688
rect 27252 68740 27304 68746
rect 27252 68682 27304 68688
rect 24872 68474 24900 68682
rect 27160 68672 27212 68678
rect 27160 68614 27212 68620
rect 23296 68468 23348 68474
rect 23296 68410 23348 68416
rect 24860 68468 24912 68474
rect 24860 68410 24912 68416
rect 23112 65408 23164 65414
rect 23112 65350 23164 65356
rect 23124 62898 23152 65350
rect 23112 62892 23164 62898
rect 23112 62834 23164 62840
rect 23308 62778 23336 68410
rect 27172 68338 27200 68614
rect 27264 68474 27292 68682
rect 27252 68468 27304 68474
rect 27252 68410 27304 68416
rect 24676 68332 24728 68338
rect 24676 68274 24728 68280
rect 27160 68332 27212 68338
rect 27160 68274 27212 68280
rect 24688 67794 24716 68274
rect 29184 68128 29236 68134
rect 29184 68070 29236 68076
rect 24676 67788 24728 67794
rect 24676 67730 24728 67736
rect 25136 66156 25188 66162
rect 25136 66098 25188 66104
rect 24400 63368 24452 63374
rect 24400 63310 24452 63316
rect 24412 62898 24440 63310
rect 24860 63300 24912 63306
rect 24860 63242 24912 63248
rect 24872 62966 24900 63242
rect 24860 62960 24912 62966
rect 24860 62902 24912 62908
rect 23388 62892 23440 62898
rect 23388 62834 23440 62840
rect 24400 62892 24452 62898
rect 24400 62834 24452 62840
rect 23124 62750 23336 62778
rect 23400 62778 23428 62834
rect 23848 62824 23900 62830
rect 23400 62750 23520 62778
rect 23848 62766 23900 62772
rect 23124 62490 23152 62750
rect 23112 62484 23164 62490
rect 23112 62426 23164 62432
rect 23124 62354 23152 62426
rect 23112 62348 23164 62354
rect 23112 62290 23164 62296
rect 22744 61736 22796 61742
rect 22744 61678 22796 61684
rect 22376 60512 22428 60518
rect 22376 60454 22428 60460
rect 22388 59634 22416 60454
rect 22376 59628 22428 59634
rect 22376 59570 22428 59576
rect 22192 59492 22244 59498
rect 22192 59434 22244 59440
rect 22204 56846 22232 59434
rect 22756 58018 22784 61678
rect 22836 60512 22888 60518
rect 22836 60454 22888 60460
rect 22848 59634 22876 60454
rect 22836 59628 22888 59634
rect 22836 59570 22888 59576
rect 22756 57990 22876 58018
rect 22468 57928 22520 57934
rect 22468 57870 22520 57876
rect 22480 57594 22508 57870
rect 22744 57860 22796 57866
rect 22744 57802 22796 57808
rect 22468 57588 22520 57594
rect 22468 57530 22520 57536
rect 22756 57526 22784 57802
rect 22744 57520 22796 57526
rect 22744 57462 22796 57468
rect 22376 57248 22428 57254
rect 22376 57190 22428 57196
rect 22192 56840 22244 56846
rect 22192 56782 22244 56788
rect 22192 56704 22244 56710
rect 22192 56646 22244 56652
rect 22204 56370 22232 56646
rect 22388 56370 22416 57190
rect 22192 56364 22244 56370
rect 22376 56364 22428 56370
rect 22244 56324 22324 56352
rect 22192 56306 22244 56312
rect 22192 55684 22244 55690
rect 22192 55626 22244 55632
rect 22204 54874 22232 55626
rect 22192 54868 22244 54874
rect 22192 54810 22244 54816
rect 22296 54534 22324 56324
rect 22376 56306 22428 56312
rect 22744 56160 22796 56166
rect 22744 56102 22796 56108
rect 22284 54528 22336 54534
rect 22284 54470 22336 54476
rect 22192 54256 22244 54262
rect 22296 54244 22324 54470
rect 22244 54216 22324 54244
rect 22192 54198 22244 54204
rect 22204 53650 22232 54198
rect 22192 53644 22244 53650
rect 22192 53586 22244 53592
rect 22204 53514 22232 53586
rect 22192 53508 22244 53514
rect 22192 53450 22244 53456
rect 22560 53508 22612 53514
rect 22560 53450 22612 53456
rect 22572 53038 22600 53450
rect 22376 53032 22428 53038
rect 22376 52974 22428 52980
rect 22560 53032 22612 53038
rect 22560 52974 22612 52980
rect 22192 51808 22244 51814
rect 22192 51750 22244 51756
rect 22204 49230 22232 51750
rect 22388 51074 22416 52974
rect 22756 52902 22784 56102
rect 22848 55962 22876 57990
rect 23020 57792 23072 57798
rect 23020 57734 23072 57740
rect 23032 57458 23060 57734
rect 23020 57452 23072 57458
rect 23020 57394 23072 57400
rect 22836 55956 22888 55962
rect 22836 55898 22888 55904
rect 22848 54806 22876 55898
rect 22928 55276 22980 55282
rect 22928 55218 22980 55224
rect 22836 54800 22888 54806
rect 22836 54742 22888 54748
rect 22836 54664 22888 54670
rect 22836 54606 22888 54612
rect 22848 53990 22876 54606
rect 22836 53984 22888 53990
rect 22836 53926 22888 53932
rect 22940 53242 22968 55218
rect 23020 54596 23072 54602
rect 23020 54538 23072 54544
rect 22928 53236 22980 53242
rect 22928 53178 22980 53184
rect 22744 52896 22796 52902
rect 22744 52838 22796 52844
rect 22468 52488 22520 52494
rect 22468 52430 22520 52436
rect 22480 51814 22508 52430
rect 22560 52420 22612 52426
rect 22560 52362 22612 52368
rect 22572 51814 22600 52362
rect 22468 51808 22520 51814
rect 22468 51750 22520 51756
rect 22560 51808 22612 51814
rect 22560 51750 22612 51756
rect 22928 51808 22980 51814
rect 22928 51750 22980 51756
rect 22388 51046 22508 51074
rect 22284 50244 22336 50250
rect 22284 50186 22336 50192
rect 22296 49910 22324 50186
rect 22376 50176 22428 50182
rect 22376 50118 22428 50124
rect 22284 49904 22336 49910
rect 22284 49846 22336 49852
rect 22192 49224 22244 49230
rect 22192 49166 22244 49172
rect 22388 49162 22416 50118
rect 22376 49156 22428 49162
rect 22376 49098 22428 49104
rect 22100 46708 22152 46714
rect 22100 46650 22152 46656
rect 22284 46572 22336 46578
rect 22284 46514 22336 46520
rect 21916 46368 21968 46374
rect 21916 46310 21968 46316
rect 21928 45966 21956 46310
rect 21916 45960 21968 45966
rect 21916 45902 21968 45908
rect 22296 45626 22324 46514
rect 22284 45620 22336 45626
rect 22284 45562 22336 45568
rect 22480 45554 22508 51046
rect 22560 50312 22612 50318
rect 22560 50254 22612 50260
rect 22572 49706 22600 50254
rect 22836 49768 22888 49774
rect 22836 49710 22888 49716
rect 22560 49700 22612 49706
rect 22560 49642 22612 49648
rect 22480 45526 22600 45554
rect 21824 44872 21876 44878
rect 21824 44814 21876 44820
rect 21836 44402 21864 44814
rect 21916 44736 21968 44742
rect 21916 44678 21968 44684
rect 21928 44470 21956 44678
rect 21916 44464 21968 44470
rect 21916 44406 21968 44412
rect 21824 44396 21876 44402
rect 21824 44338 21876 44344
rect 21836 43790 21864 44338
rect 21824 43784 21876 43790
rect 21824 43726 21876 43732
rect 21928 43722 21956 44406
rect 22008 44192 22060 44198
rect 22008 44134 22060 44140
rect 21916 43716 21968 43722
rect 21916 43658 21968 43664
rect 21824 41540 21876 41546
rect 21824 41482 21876 41488
rect 21836 41274 21864 41482
rect 21916 41472 21968 41478
rect 21916 41414 21968 41420
rect 21824 41268 21876 41274
rect 21824 41210 21876 41216
rect 21928 41070 21956 41414
rect 21916 41064 21968 41070
rect 21916 41006 21968 41012
rect 22020 40662 22048 44134
rect 22572 43314 22600 45526
rect 22744 43784 22796 43790
rect 22744 43726 22796 43732
rect 22560 43308 22612 43314
rect 22560 43250 22612 43256
rect 22756 42906 22784 43726
rect 22744 42900 22796 42906
rect 22744 42842 22796 42848
rect 22284 42628 22336 42634
rect 22284 42570 22336 42576
rect 22100 42152 22152 42158
rect 22100 42094 22152 42100
rect 22112 41682 22140 42094
rect 22100 41676 22152 41682
rect 22100 41618 22152 41624
rect 22296 41138 22324 42570
rect 22466 41576 22522 41585
rect 22466 41511 22522 41520
rect 22284 41132 22336 41138
rect 22192 41116 22244 41122
rect 22284 41074 22336 41080
rect 22192 41058 22244 41064
rect 22204 40730 22232 41058
rect 22192 40724 22244 40730
rect 22192 40666 22244 40672
rect 22008 40656 22060 40662
rect 22008 40598 22060 40604
rect 22480 40186 22508 41511
rect 22744 40724 22796 40730
rect 22744 40666 22796 40672
rect 22468 40180 22520 40186
rect 22468 40122 22520 40128
rect 22480 39506 22508 40122
rect 22468 39500 22520 39506
rect 22388 39460 22468 39488
rect 22388 38350 22416 39460
rect 22468 39442 22520 39448
rect 22560 39364 22612 39370
rect 22560 39306 22612 39312
rect 22572 39098 22600 39306
rect 22560 39092 22612 39098
rect 22560 39034 22612 39040
rect 22756 38894 22784 40666
rect 22848 40050 22876 49710
rect 22836 40044 22888 40050
rect 22836 39986 22888 39992
rect 22744 38888 22796 38894
rect 22744 38830 22796 38836
rect 22376 38344 22428 38350
rect 22376 38286 22428 38292
rect 22744 37188 22796 37194
rect 22744 37130 22796 37136
rect 22756 36922 22784 37130
rect 22940 37126 22968 51750
rect 23032 50318 23060 54538
rect 23124 50980 23152 62290
rect 23204 57452 23256 57458
rect 23204 57394 23256 57400
rect 23216 57050 23244 57394
rect 23204 57044 23256 57050
rect 23204 56986 23256 56992
rect 23204 55752 23256 55758
rect 23204 55694 23256 55700
rect 23216 54194 23244 55694
rect 23388 54664 23440 54670
rect 23388 54606 23440 54612
rect 23296 54528 23348 54534
rect 23296 54470 23348 54476
rect 23308 54194 23336 54470
rect 23204 54188 23256 54194
rect 23204 54130 23256 54136
rect 23296 54188 23348 54194
rect 23296 54130 23348 54136
rect 23216 52494 23244 54130
rect 23400 53786 23428 54606
rect 23388 53780 23440 53786
rect 23388 53722 23440 53728
rect 23296 53236 23348 53242
rect 23296 53178 23348 53184
rect 23204 52488 23256 52494
rect 23204 52430 23256 52436
rect 23124 50952 23244 50980
rect 23020 50312 23072 50318
rect 23020 50254 23072 50260
rect 23020 49700 23072 49706
rect 23020 49642 23072 49648
rect 23032 49434 23060 49642
rect 23020 49428 23072 49434
rect 23020 49370 23072 49376
rect 23112 47660 23164 47666
rect 23112 47602 23164 47608
rect 23124 47258 23152 47602
rect 23112 47252 23164 47258
rect 23112 47194 23164 47200
rect 23020 43648 23072 43654
rect 23020 43590 23072 43596
rect 23032 38962 23060 43590
rect 23112 41472 23164 41478
rect 23112 41414 23164 41420
rect 23124 39098 23152 41414
rect 23112 39092 23164 39098
rect 23112 39034 23164 39040
rect 23020 38956 23072 38962
rect 23020 38898 23072 38904
rect 23124 38894 23152 39034
rect 23112 38888 23164 38894
rect 23112 38830 23164 38836
rect 22928 37120 22980 37126
rect 22928 37062 22980 37068
rect 22744 36916 22796 36922
rect 22744 36858 22796 36864
rect 22284 36168 22336 36174
rect 22284 36110 22336 36116
rect 22296 35290 22324 36110
rect 23020 36100 23072 36106
rect 23020 36042 23072 36048
rect 22652 35692 22704 35698
rect 22652 35634 22704 35640
rect 22560 35624 22612 35630
rect 22560 35566 22612 35572
rect 21732 35284 21784 35290
rect 21732 35226 21784 35232
rect 22284 35284 22336 35290
rect 22284 35226 22336 35232
rect 22376 35080 22428 35086
rect 22376 35022 22428 35028
rect 22388 33522 22416 35022
rect 22468 33992 22520 33998
rect 22468 33934 22520 33940
rect 22480 33658 22508 33934
rect 22468 33652 22520 33658
rect 22468 33594 22520 33600
rect 22376 33516 22428 33522
rect 22376 33458 22428 33464
rect 22388 32994 22416 33458
rect 22388 32966 22508 32994
rect 22376 32360 22428 32366
rect 22376 32302 22428 32308
rect 22388 32026 22416 32302
rect 22376 32020 22428 32026
rect 22376 31962 22428 31968
rect 22480 31822 22508 32966
rect 22468 31816 22520 31822
rect 22468 31758 22520 31764
rect 22480 31482 22508 31758
rect 22468 31476 22520 31482
rect 22468 31418 22520 31424
rect 22468 30728 22520 30734
rect 22468 30670 22520 30676
rect 22100 30592 22152 30598
rect 22100 30534 22152 30540
rect 21824 30048 21876 30054
rect 21824 29990 21876 29996
rect 21836 29714 21864 29990
rect 21824 29708 21876 29714
rect 21824 29650 21876 29656
rect 22112 29646 22140 30534
rect 22480 30394 22508 30670
rect 22468 30388 22520 30394
rect 22468 30330 22520 30336
rect 22100 29640 22152 29646
rect 22100 29582 22152 29588
rect 22572 12646 22600 35566
rect 22664 35222 22692 35634
rect 23032 35290 23060 36042
rect 23020 35284 23072 35290
rect 23020 35226 23072 35232
rect 22652 35216 22704 35222
rect 22652 35158 22704 35164
rect 22744 34400 22796 34406
rect 22744 34342 22796 34348
rect 22756 33998 22784 34342
rect 22744 33992 22796 33998
rect 22744 33934 22796 33940
rect 22836 32768 22888 32774
rect 22836 32710 22888 32716
rect 22848 32502 22876 32710
rect 22836 32496 22888 32502
rect 22836 32438 22888 32444
rect 23020 32224 23072 32230
rect 23020 32166 23072 32172
rect 23032 31890 23060 32166
rect 23020 31884 23072 31890
rect 23020 31826 23072 31832
rect 23216 31754 23244 50952
rect 23308 49230 23336 53178
rect 23492 50318 23520 62750
rect 23572 61736 23624 61742
rect 23572 61678 23624 61684
rect 23584 61402 23612 61678
rect 23572 61396 23624 61402
rect 23572 61338 23624 61344
rect 23664 60580 23716 60586
rect 23664 60522 23716 60528
rect 23676 57458 23704 60522
rect 23756 60104 23808 60110
rect 23756 60046 23808 60052
rect 23664 57452 23716 57458
rect 23664 57394 23716 57400
rect 23676 52630 23704 57394
rect 23664 52624 23716 52630
rect 23664 52566 23716 52572
rect 23664 52420 23716 52426
rect 23664 52362 23716 52368
rect 23676 52086 23704 52362
rect 23664 52080 23716 52086
rect 23664 52022 23716 52028
rect 23768 51066 23796 60046
rect 23756 51060 23808 51066
rect 23756 51002 23808 51008
rect 23388 50312 23440 50318
rect 23388 50254 23440 50260
rect 23480 50312 23532 50318
rect 23480 50254 23532 50260
rect 23296 49224 23348 49230
rect 23296 49166 23348 49172
rect 23296 49088 23348 49094
rect 23296 49030 23348 49036
rect 23308 48142 23336 49030
rect 23296 48136 23348 48142
rect 23296 48078 23348 48084
rect 23296 48000 23348 48006
rect 23296 47942 23348 47948
rect 23308 47054 23336 47942
rect 23296 47048 23348 47054
rect 23296 46990 23348 46996
rect 23296 45416 23348 45422
rect 23296 45358 23348 45364
rect 23308 44538 23336 45358
rect 23296 44532 23348 44538
rect 23296 44474 23348 44480
rect 23400 42226 23428 50254
rect 23388 42220 23440 42226
rect 23388 42162 23440 42168
rect 23400 41478 23428 42162
rect 23388 41472 23440 41478
rect 23388 41414 23440 41420
rect 23296 41268 23348 41274
rect 23296 41210 23348 41216
rect 23308 40526 23336 41210
rect 23492 41206 23520 50254
rect 23664 48068 23716 48074
rect 23664 48010 23716 48016
rect 23676 47462 23704 48010
rect 23664 47456 23716 47462
rect 23664 47398 23716 47404
rect 23664 45824 23716 45830
rect 23664 45766 23716 45772
rect 23676 45558 23704 45766
rect 23664 45552 23716 45558
rect 23664 45494 23716 45500
rect 23572 44872 23624 44878
rect 23572 44814 23624 44820
rect 23584 44402 23612 44814
rect 23572 44396 23624 44402
rect 23572 44338 23624 44344
rect 23664 42560 23716 42566
rect 23664 42502 23716 42508
rect 23572 42152 23624 42158
rect 23572 42094 23624 42100
rect 23584 41614 23612 42094
rect 23676 41818 23704 42502
rect 23664 41812 23716 41818
rect 23664 41754 23716 41760
rect 23572 41608 23624 41614
rect 23572 41550 23624 41556
rect 23480 41200 23532 41206
rect 23480 41142 23532 41148
rect 23676 41138 23704 41754
rect 23664 41132 23716 41138
rect 23664 41074 23716 41080
rect 23676 40594 23704 41074
rect 23664 40588 23716 40594
rect 23664 40530 23716 40536
rect 23296 40520 23348 40526
rect 23296 40462 23348 40468
rect 23308 37874 23336 40462
rect 23388 40384 23440 40390
rect 23388 40326 23440 40332
rect 23400 40118 23428 40326
rect 23388 40112 23440 40118
rect 23388 40054 23440 40060
rect 23400 38350 23428 40054
rect 23756 39296 23808 39302
rect 23756 39238 23808 39244
rect 23768 38962 23796 39238
rect 23756 38956 23808 38962
rect 23756 38898 23808 38904
rect 23388 38344 23440 38350
rect 23388 38286 23440 38292
rect 23296 37868 23348 37874
rect 23296 37810 23348 37816
rect 23308 36786 23336 37810
rect 23296 36780 23348 36786
rect 23296 36722 23348 36728
rect 23572 36168 23624 36174
rect 23572 36110 23624 36116
rect 23480 34604 23532 34610
rect 23480 34546 23532 34552
rect 23388 34196 23440 34202
rect 23388 34138 23440 34144
rect 23400 33590 23428 34138
rect 23492 33658 23520 34546
rect 23480 33652 23532 33658
rect 23480 33594 23532 33600
rect 23388 33584 23440 33590
rect 23388 33526 23440 33532
rect 23584 33522 23612 36110
rect 23756 36032 23808 36038
rect 23756 35974 23808 35980
rect 23768 35086 23796 35974
rect 23756 35080 23808 35086
rect 23756 35022 23808 35028
rect 23572 33516 23624 33522
rect 23572 33458 23624 33464
rect 23388 32904 23440 32910
rect 23388 32846 23440 32852
rect 23400 32026 23428 32846
rect 23388 32020 23440 32026
rect 23388 31962 23440 31968
rect 23584 31890 23612 33458
rect 23572 31884 23624 31890
rect 23572 31826 23624 31832
rect 23124 31726 23244 31754
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 23124 3602 23152 31726
rect 23204 31476 23256 31482
rect 23204 31418 23256 31424
rect 23216 30734 23244 31418
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23216 30326 23244 30670
rect 23480 30660 23532 30666
rect 23480 30602 23532 30608
rect 23204 30320 23256 30326
rect 23204 30262 23256 30268
rect 23492 30258 23520 30602
rect 23584 30326 23612 31826
rect 23572 30320 23624 30326
rect 23572 30262 23624 30268
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 23204 30184 23256 30190
rect 23204 30126 23256 30132
rect 23216 29850 23244 30126
rect 23204 29844 23256 29850
rect 23204 29786 23256 29792
rect 23584 29646 23612 30262
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 23204 28008 23256 28014
rect 23204 27950 23256 27956
rect 23216 27674 23244 27950
rect 23204 27668 23256 27674
rect 23204 27610 23256 27616
rect 23112 3596 23164 3602
rect 23112 3538 23164 3544
rect 23860 3534 23888 62766
rect 24412 62286 24440 62834
rect 24400 62280 24452 62286
rect 24400 62222 24452 62228
rect 24308 61600 24360 61606
rect 24308 61542 24360 61548
rect 24320 58546 24348 61542
rect 24412 61198 24440 62222
rect 24872 61266 24900 62902
rect 25148 61878 25176 66098
rect 25320 63504 25372 63510
rect 25320 63446 25372 63452
rect 25332 62218 25360 63446
rect 29092 62824 29144 62830
rect 29196 62812 29224 68070
rect 29276 62824 29328 62830
rect 29196 62784 29276 62812
rect 29092 62766 29144 62772
rect 29276 62766 29328 62772
rect 26240 62280 26292 62286
rect 26240 62222 26292 62228
rect 29000 62280 29052 62286
rect 29000 62222 29052 62228
rect 25320 62212 25372 62218
rect 25320 62154 25372 62160
rect 25964 62212 26016 62218
rect 25964 62154 26016 62160
rect 25136 61872 25188 61878
rect 25136 61814 25188 61820
rect 24860 61260 24912 61266
rect 24860 61202 24912 61208
rect 24400 61192 24452 61198
rect 24400 61134 24452 61140
rect 24952 60512 25004 60518
rect 24952 60454 25004 60460
rect 24964 60110 24992 60454
rect 24952 60104 25004 60110
rect 24952 60046 25004 60052
rect 25228 58880 25280 58886
rect 25228 58822 25280 58828
rect 24308 58540 24360 58546
rect 24308 58482 24360 58488
rect 24584 58336 24636 58342
rect 24584 58278 24636 58284
rect 24596 58002 24624 58278
rect 24584 57996 24636 58002
rect 24584 57938 24636 57944
rect 25240 57526 25268 58822
rect 25228 57520 25280 57526
rect 25228 57462 25280 57468
rect 24952 57452 25004 57458
rect 24952 57394 25004 57400
rect 24216 57384 24268 57390
rect 24216 57326 24268 57332
rect 24228 57050 24256 57326
rect 24216 57044 24268 57050
rect 24216 56986 24268 56992
rect 24964 56370 24992 57394
rect 25044 56772 25096 56778
rect 25044 56714 25096 56720
rect 24952 56364 25004 56370
rect 24952 56306 25004 56312
rect 24492 56160 24544 56166
rect 24492 56102 24544 56108
rect 24504 55826 24532 56102
rect 24492 55820 24544 55826
rect 24492 55762 24544 55768
rect 24032 54732 24084 54738
rect 24032 54674 24084 54680
rect 24044 52970 24072 54674
rect 24964 54194 24992 56306
rect 24952 54188 25004 54194
rect 24952 54130 25004 54136
rect 24860 53984 24912 53990
rect 24860 53926 24912 53932
rect 24872 53650 24900 53926
rect 24860 53644 24912 53650
rect 24860 53586 24912 53592
rect 24860 53168 24912 53174
rect 24860 53110 24912 53116
rect 24400 53100 24452 53106
rect 24400 53042 24452 53048
rect 24032 52964 24084 52970
rect 24032 52906 24084 52912
rect 24044 51882 24072 52906
rect 24412 52698 24440 53042
rect 24492 52964 24544 52970
rect 24492 52906 24544 52912
rect 24400 52692 24452 52698
rect 24400 52634 24452 52640
rect 24308 52624 24360 52630
rect 24308 52566 24360 52572
rect 24216 52488 24268 52494
rect 24216 52430 24268 52436
rect 24124 52352 24176 52358
rect 24124 52294 24176 52300
rect 24032 51876 24084 51882
rect 24032 51818 24084 51824
rect 24044 51066 24072 51818
rect 24136 51814 24164 52294
rect 24124 51808 24176 51814
rect 24124 51750 24176 51756
rect 24032 51060 24084 51066
rect 24032 51002 24084 51008
rect 24044 50318 24072 51002
rect 24136 50386 24164 51750
rect 24124 50380 24176 50386
rect 24124 50322 24176 50328
rect 24032 50312 24084 50318
rect 24032 50254 24084 50260
rect 24032 46912 24084 46918
rect 24032 46854 24084 46860
rect 24044 46578 24072 46854
rect 24032 46572 24084 46578
rect 24032 46514 24084 46520
rect 24032 46164 24084 46170
rect 24032 46106 24084 46112
rect 24044 44470 24072 46106
rect 24032 44464 24084 44470
rect 24032 44406 24084 44412
rect 24032 44328 24084 44334
rect 24032 44270 24084 44276
rect 24044 43314 24072 44270
rect 24124 43784 24176 43790
rect 24124 43726 24176 43732
rect 24136 43450 24164 43726
rect 24124 43444 24176 43450
rect 24124 43386 24176 43392
rect 24032 43308 24084 43314
rect 24032 43250 24084 43256
rect 24044 42634 24072 43250
rect 24032 42628 24084 42634
rect 24032 42570 24084 42576
rect 24044 42022 24072 42570
rect 24228 42158 24256 52430
rect 24320 52018 24348 52566
rect 24308 52012 24360 52018
rect 24308 51954 24360 51960
rect 24412 51270 24440 52634
rect 24504 52494 24532 52906
rect 24584 52896 24636 52902
rect 24584 52838 24636 52844
rect 24492 52488 24544 52494
rect 24492 52430 24544 52436
rect 24596 51950 24624 52838
rect 24872 52018 24900 53110
rect 24860 52012 24912 52018
rect 24860 51954 24912 51960
rect 24584 51944 24636 51950
rect 24584 51886 24636 51892
rect 24768 51808 24820 51814
rect 24768 51750 24820 51756
rect 24780 51474 24808 51750
rect 24768 51468 24820 51474
rect 24768 51410 24820 51416
rect 24964 51338 24992 54130
rect 24952 51332 25004 51338
rect 24952 51274 25004 51280
rect 24400 51264 24452 51270
rect 24400 51206 24452 51212
rect 24400 50924 24452 50930
rect 24400 50866 24452 50872
rect 24676 50924 24728 50930
rect 24676 50866 24728 50872
rect 24412 50522 24440 50866
rect 24400 50516 24452 50522
rect 24400 50458 24452 50464
rect 24412 49842 24440 50458
rect 24400 49836 24452 49842
rect 24400 49778 24452 49784
rect 24308 48136 24360 48142
rect 24308 48078 24360 48084
rect 24320 47802 24348 48078
rect 24308 47796 24360 47802
rect 24308 47738 24360 47744
rect 24308 47660 24360 47666
rect 24308 47602 24360 47608
rect 24320 43654 24348 47602
rect 24688 46322 24716 50866
rect 24964 49978 24992 51274
rect 25056 50930 25084 56714
rect 25332 56250 25360 62154
rect 25976 61810 26004 62154
rect 26252 61946 26280 62222
rect 26516 62212 26568 62218
rect 26516 62154 26568 62160
rect 26240 61940 26292 61946
rect 26240 61882 26292 61888
rect 26056 61872 26108 61878
rect 26056 61814 26108 61820
rect 25688 61804 25740 61810
rect 25688 61746 25740 61752
rect 25964 61804 26016 61810
rect 25964 61746 26016 61752
rect 25504 60716 25556 60722
rect 25504 60658 25556 60664
rect 25516 59770 25544 60658
rect 25504 59764 25556 59770
rect 25504 59706 25556 59712
rect 25412 59628 25464 59634
rect 25412 59570 25464 59576
rect 25424 58546 25452 59570
rect 25596 59016 25648 59022
rect 25596 58958 25648 58964
rect 25608 58682 25636 58958
rect 25596 58676 25648 58682
rect 25596 58618 25648 58624
rect 25412 58540 25464 58546
rect 25412 58482 25464 58488
rect 25424 56522 25452 58482
rect 25424 56494 25544 56522
rect 25412 56364 25464 56370
rect 25412 56306 25464 56312
rect 25240 56222 25360 56250
rect 25136 55616 25188 55622
rect 25136 55558 25188 55564
rect 25148 55282 25176 55558
rect 25136 55276 25188 55282
rect 25136 55218 25188 55224
rect 25136 54528 25188 54534
rect 25136 54470 25188 54476
rect 25148 53582 25176 54470
rect 25136 53576 25188 53582
rect 25136 53518 25188 53524
rect 25136 52352 25188 52358
rect 25136 52294 25188 52300
rect 25148 51406 25176 52294
rect 25136 51400 25188 51406
rect 25136 51342 25188 51348
rect 25044 50924 25096 50930
rect 25044 50866 25096 50872
rect 24952 49972 25004 49978
rect 24952 49914 25004 49920
rect 25136 49972 25188 49978
rect 25136 49914 25188 49920
rect 24860 49224 24912 49230
rect 24964 49212 24992 49914
rect 24912 49184 24992 49212
rect 24860 49166 24912 49172
rect 24860 48680 24912 48686
rect 24860 48622 24912 48628
rect 24872 48006 24900 48622
rect 24860 48000 24912 48006
rect 24860 47942 24912 47948
rect 24768 47456 24820 47462
rect 24768 47398 24820 47404
rect 24780 46594 24808 47398
rect 24872 46918 24900 47942
rect 24860 46912 24912 46918
rect 24860 46854 24912 46860
rect 24780 46578 24992 46594
rect 24780 46572 25004 46578
rect 24780 46566 24952 46572
rect 24952 46514 25004 46520
rect 24768 46504 24820 46510
rect 25044 46504 25096 46510
rect 24820 46452 24900 46458
rect 24768 46446 24900 46452
rect 25044 46446 25096 46452
rect 24780 46430 24900 46446
rect 24688 46294 24808 46322
rect 24676 45892 24728 45898
rect 24676 45834 24728 45840
rect 24688 45626 24716 45834
rect 24780 45626 24808 46294
rect 24676 45620 24728 45626
rect 24676 45562 24728 45568
rect 24768 45620 24820 45626
rect 24768 45562 24820 45568
rect 24872 45558 24900 46430
rect 24952 45960 25004 45966
rect 24952 45902 25004 45908
rect 24964 45778 24992 45902
rect 25056 45898 25084 46446
rect 25044 45892 25096 45898
rect 25044 45834 25096 45840
rect 25148 45778 25176 49914
rect 24964 45750 25176 45778
rect 24860 45552 24912 45558
rect 25240 45554 25268 56222
rect 25320 56160 25372 56166
rect 25320 56102 25372 56108
rect 25332 55758 25360 56102
rect 25320 55752 25372 55758
rect 25320 55694 25372 55700
rect 25424 55418 25452 56306
rect 25412 55412 25464 55418
rect 25412 55354 25464 55360
rect 25516 55282 25544 56494
rect 25700 55282 25728 61746
rect 25872 61736 25924 61742
rect 25872 61678 25924 61684
rect 25884 61130 25912 61678
rect 25872 61124 25924 61130
rect 25872 61066 25924 61072
rect 25884 60734 25912 61066
rect 25884 60706 26004 60734
rect 25780 60308 25832 60314
rect 25780 60250 25832 60256
rect 25792 59702 25820 60250
rect 25780 59696 25832 59702
rect 25780 59638 25832 59644
rect 25504 55276 25556 55282
rect 25504 55218 25556 55224
rect 25688 55276 25740 55282
rect 25688 55218 25740 55224
rect 25412 54664 25464 54670
rect 25412 54606 25464 54612
rect 25424 53242 25452 54606
rect 25412 53236 25464 53242
rect 25412 53178 25464 53184
rect 25516 53106 25544 55218
rect 25504 53100 25556 53106
rect 25504 53042 25556 53048
rect 25412 52488 25464 52494
rect 25412 52430 25464 52436
rect 25320 52012 25372 52018
rect 25320 51954 25372 51960
rect 25332 50862 25360 51954
rect 25424 51066 25452 52430
rect 25516 52018 25544 53042
rect 25504 52012 25556 52018
rect 25504 51954 25556 51960
rect 25504 51876 25556 51882
rect 25504 51818 25556 51824
rect 25412 51060 25464 51066
rect 25412 51002 25464 51008
rect 25320 50856 25372 50862
rect 25320 50798 25372 50804
rect 25516 49978 25544 51818
rect 25872 50244 25924 50250
rect 25872 50186 25924 50192
rect 25504 49972 25556 49978
rect 25504 49914 25556 49920
rect 25884 49745 25912 50186
rect 25870 49736 25926 49745
rect 25870 49671 25926 49680
rect 25412 48544 25464 48550
rect 25412 48486 25464 48492
rect 25424 48142 25452 48486
rect 25412 48136 25464 48142
rect 25412 48078 25464 48084
rect 25872 48000 25924 48006
rect 25872 47942 25924 47948
rect 25884 47734 25912 47942
rect 25872 47728 25924 47734
rect 25872 47670 25924 47676
rect 25872 47592 25924 47598
rect 25872 47534 25924 47540
rect 25596 46980 25648 46986
rect 25596 46922 25648 46928
rect 25608 46050 25636 46922
rect 25688 46368 25740 46374
rect 25688 46310 25740 46316
rect 25700 46170 25728 46310
rect 25688 46164 25740 46170
rect 25688 46106 25740 46112
rect 25608 46022 25728 46050
rect 25504 45892 25556 45898
rect 25504 45834 25556 45840
rect 25240 45526 25360 45554
rect 24860 45494 24912 45500
rect 25228 44396 25280 44402
rect 25228 44338 25280 44344
rect 25044 44192 25096 44198
rect 25044 44134 25096 44140
rect 25056 43790 25084 44134
rect 25044 43784 25096 43790
rect 25044 43726 25096 43732
rect 24308 43648 24360 43654
rect 24308 43590 24360 43596
rect 24216 42152 24268 42158
rect 24216 42094 24268 42100
rect 24320 42090 24348 43590
rect 25240 43450 25268 44338
rect 25228 43444 25280 43450
rect 25228 43386 25280 43392
rect 25228 43240 25280 43246
rect 25228 43182 25280 43188
rect 25044 42696 25096 42702
rect 25044 42638 25096 42644
rect 24492 42628 24544 42634
rect 24492 42570 24544 42576
rect 24308 42084 24360 42090
rect 24308 42026 24360 42032
rect 24032 42016 24084 42022
rect 24032 41958 24084 41964
rect 24044 41206 24072 41958
rect 24504 41818 24532 42570
rect 24952 42560 25004 42566
rect 24952 42502 25004 42508
rect 24964 42226 24992 42502
rect 25056 42362 25084 42638
rect 25044 42356 25096 42362
rect 25044 42298 25096 42304
rect 25240 42226 25268 43182
rect 24952 42220 25004 42226
rect 24952 42162 25004 42168
rect 25228 42220 25280 42226
rect 25228 42162 25280 42168
rect 24584 42016 24636 42022
rect 24584 41958 24636 41964
rect 24492 41812 24544 41818
rect 24492 41754 24544 41760
rect 24596 41614 24624 41958
rect 24584 41608 24636 41614
rect 24584 41550 24636 41556
rect 24032 41200 24084 41206
rect 24032 41142 24084 41148
rect 24952 41132 25004 41138
rect 24952 41074 25004 41080
rect 24400 40996 24452 41002
rect 24400 40938 24452 40944
rect 24412 40594 24440 40938
rect 24676 40928 24728 40934
rect 24676 40870 24728 40876
rect 24400 40588 24452 40594
rect 24400 40530 24452 40536
rect 24688 40526 24716 40870
rect 24676 40520 24728 40526
rect 24676 40462 24728 40468
rect 24964 40186 24992 41074
rect 25136 40384 25188 40390
rect 25136 40326 25188 40332
rect 24952 40180 25004 40186
rect 24952 40122 25004 40128
rect 25148 40050 25176 40326
rect 25240 40050 25268 42162
rect 25136 40044 25188 40050
rect 25136 39986 25188 39992
rect 25228 40044 25280 40050
rect 25228 39986 25280 39992
rect 25240 39030 25268 39986
rect 25228 39024 25280 39030
rect 25228 38966 25280 38972
rect 24032 38888 24084 38894
rect 24032 38830 24084 38836
rect 24044 38554 24072 38830
rect 24032 38548 24084 38554
rect 24032 38490 24084 38496
rect 24400 38344 24452 38350
rect 24400 38286 24452 38292
rect 24412 38010 24440 38286
rect 24676 38276 24728 38282
rect 24676 38218 24728 38224
rect 24400 38004 24452 38010
rect 24400 37946 24452 37952
rect 24216 37800 24268 37806
rect 24216 37742 24268 37748
rect 24228 26790 24256 37742
rect 24688 36922 24716 38218
rect 25332 37754 25360 45526
rect 25516 45082 25544 45834
rect 25596 45824 25648 45830
rect 25596 45766 25648 45772
rect 25608 45558 25636 45766
rect 25700 45558 25728 46022
rect 25780 45960 25832 45966
rect 25780 45902 25832 45908
rect 25596 45552 25648 45558
rect 25596 45494 25648 45500
rect 25688 45552 25740 45558
rect 25688 45494 25740 45500
rect 25792 45422 25820 45902
rect 25780 45416 25832 45422
rect 25780 45358 25832 45364
rect 25504 45076 25556 45082
rect 25504 45018 25556 45024
rect 25412 43920 25464 43926
rect 25412 43862 25464 43868
rect 25424 43314 25452 43862
rect 25780 43376 25832 43382
rect 25780 43318 25832 43324
rect 25412 43308 25464 43314
rect 25412 43250 25464 43256
rect 25688 42764 25740 42770
rect 25688 42706 25740 42712
rect 25412 42220 25464 42226
rect 25412 42162 25464 42168
rect 25240 37726 25360 37754
rect 24860 37120 24912 37126
rect 24860 37062 24912 37068
rect 24676 36916 24728 36922
rect 24676 36858 24728 36864
rect 24872 36786 24900 37062
rect 24860 36780 24912 36786
rect 24860 36722 24912 36728
rect 24308 36576 24360 36582
rect 24308 36518 24360 36524
rect 24320 27470 24348 36518
rect 24492 35692 24544 35698
rect 24492 35634 24544 35640
rect 24504 34746 24532 35634
rect 24860 34944 24912 34950
rect 24860 34886 24912 34892
rect 24492 34740 24544 34746
rect 24492 34682 24544 34688
rect 24872 34610 24900 34886
rect 24860 34604 24912 34610
rect 24860 34546 24912 34552
rect 24952 33992 25004 33998
rect 24952 33934 25004 33940
rect 24400 33856 24452 33862
rect 24400 33798 24452 33804
rect 24412 33522 24440 33798
rect 24400 33516 24452 33522
rect 24400 33458 24452 33464
rect 24964 33114 24992 33934
rect 25136 33856 25188 33862
rect 25136 33798 25188 33804
rect 25148 33590 25176 33798
rect 25136 33584 25188 33590
rect 25136 33526 25188 33532
rect 24952 33108 25004 33114
rect 24952 33050 25004 33056
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24400 30592 24452 30598
rect 24400 30534 24452 30540
rect 24412 30326 24440 30534
rect 24400 30320 24452 30326
rect 24400 30262 24452 30268
rect 24492 30116 24544 30122
rect 24492 30058 24544 30064
rect 24400 30048 24452 30054
rect 24400 29990 24452 29996
rect 24412 29714 24440 29990
rect 24504 29850 24532 30058
rect 24596 29850 24624 30670
rect 24492 29844 24544 29850
rect 24492 29786 24544 29792
rect 24584 29844 24636 29850
rect 24584 29786 24636 29792
rect 24400 29708 24452 29714
rect 24400 29650 24452 29656
rect 24676 29096 24728 29102
rect 24676 29038 24728 29044
rect 24688 28762 24716 29038
rect 24676 28756 24728 28762
rect 24676 28698 24728 28704
rect 24964 28490 24992 33050
rect 25240 31754 25268 37726
rect 25320 37664 25372 37670
rect 25320 37606 25372 37612
rect 25332 37330 25360 37606
rect 25320 37324 25372 37330
rect 25320 37266 25372 37272
rect 25320 36032 25372 36038
rect 25320 35974 25372 35980
rect 25332 35766 25360 35974
rect 25320 35760 25372 35766
rect 25320 35702 25372 35708
rect 25320 35080 25372 35086
rect 25320 35022 25372 35028
rect 25332 34746 25360 35022
rect 25320 34740 25372 34746
rect 25320 34682 25372 34688
rect 25320 33992 25372 33998
rect 25320 33934 25372 33940
rect 25332 32570 25360 33934
rect 25320 32564 25372 32570
rect 25320 32506 25372 32512
rect 25240 31726 25360 31754
rect 25044 31680 25096 31686
rect 25044 31622 25096 31628
rect 25056 31346 25084 31622
rect 25044 31340 25096 31346
rect 25044 31282 25096 31288
rect 25228 29504 25280 29510
rect 25228 29446 25280 29452
rect 25240 29238 25268 29446
rect 25228 29232 25280 29238
rect 25228 29174 25280 29180
rect 24952 28484 25004 28490
rect 24952 28426 25004 28432
rect 24308 27464 24360 27470
rect 24308 27406 24360 27412
rect 24320 26994 24348 27406
rect 24584 27396 24636 27402
rect 24584 27338 24636 27344
rect 24596 27130 24624 27338
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24308 26988 24360 26994
rect 24308 26930 24360 26936
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 24228 26234 24256 26726
rect 24320 26518 24348 26930
rect 24308 26512 24360 26518
rect 24308 26454 24360 26460
rect 24136 26206 24256 26234
rect 24136 4622 24164 26206
rect 24124 4616 24176 4622
rect 24124 4558 24176 4564
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 22112 3126 22140 3334
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 22560 2916 22612 2922
rect 22560 2858 22612 2864
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 20904 2372 20956 2378
rect 20904 2314 20956 2320
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 21284 800 21312 2382
rect 22572 800 22600 2858
rect 22756 2650 22784 2926
rect 22744 2644 22796 2650
rect 22744 2586 22796 2592
rect 24504 800 24532 3334
rect 25332 2514 25360 31726
rect 25424 2582 25452 42162
rect 25596 38888 25648 38894
rect 25596 38830 25648 38836
rect 25504 37120 25556 37126
rect 25504 37062 25556 37068
rect 25516 36786 25544 37062
rect 25504 36780 25556 36786
rect 25504 36722 25556 36728
rect 25516 35018 25544 36722
rect 25504 35012 25556 35018
rect 25504 34954 25556 34960
rect 25516 32434 25544 34954
rect 25504 32428 25556 32434
rect 25504 32370 25556 32376
rect 25516 28558 25544 32370
rect 25504 28552 25556 28558
rect 25504 28494 25556 28500
rect 25516 28150 25544 28494
rect 25504 28144 25556 28150
rect 25504 28086 25556 28092
rect 25608 3466 25636 38830
rect 25700 36854 25728 42706
rect 25792 41818 25820 43318
rect 25884 42362 25912 47534
rect 25976 45554 26004 60706
rect 26068 51074 26096 61814
rect 26528 61402 26556 62154
rect 27436 62144 27488 62150
rect 27436 62086 27488 62092
rect 28264 62144 28316 62150
rect 28264 62086 28316 62092
rect 28816 62144 28868 62150
rect 28816 62086 28868 62092
rect 26516 61396 26568 61402
rect 26516 61338 26568 61344
rect 27448 61198 27476 62086
rect 28276 61810 28304 62086
rect 28828 61878 28856 62086
rect 28816 61872 28868 61878
rect 28816 61814 28868 61820
rect 28264 61804 28316 61810
rect 28264 61746 28316 61752
rect 27804 61600 27856 61606
rect 27804 61542 27856 61548
rect 27896 61600 27948 61606
rect 27896 61542 27948 61548
rect 27816 61334 27844 61542
rect 27804 61328 27856 61334
rect 27804 61270 27856 61276
rect 27908 61198 27936 61542
rect 29012 61402 29040 62222
rect 29000 61396 29052 61402
rect 29000 61338 29052 61344
rect 27436 61192 27488 61198
rect 27436 61134 27488 61140
rect 27896 61192 27948 61198
rect 27896 61134 27948 61140
rect 28356 61192 28408 61198
rect 28356 61134 28408 61140
rect 26240 60852 26292 60858
rect 26240 60794 26292 60800
rect 26252 59702 26280 60794
rect 26332 60648 26384 60654
rect 26332 60590 26384 60596
rect 26344 60110 26372 60590
rect 27448 60178 27476 61134
rect 27712 60716 27764 60722
rect 27712 60658 27764 60664
rect 27620 60240 27672 60246
rect 27620 60182 27672 60188
rect 27436 60172 27488 60178
rect 27436 60114 27488 60120
rect 26332 60104 26384 60110
rect 26384 60064 26464 60092
rect 26332 60046 26384 60052
rect 26332 59968 26384 59974
rect 26332 59910 26384 59916
rect 26344 59770 26372 59910
rect 26332 59764 26384 59770
rect 26332 59706 26384 59712
rect 26240 59696 26292 59702
rect 26240 59638 26292 59644
rect 26240 58676 26292 58682
rect 26240 58618 26292 58624
rect 26146 58032 26202 58041
rect 26146 57967 26148 57976
rect 26200 57967 26202 57976
rect 26148 57938 26200 57944
rect 26252 57322 26280 58618
rect 26436 58546 26464 60064
rect 26976 59968 27028 59974
rect 26976 59910 27028 59916
rect 26988 59634 27016 59910
rect 27632 59634 27660 60182
rect 26976 59628 27028 59634
rect 26976 59570 27028 59576
rect 27620 59628 27672 59634
rect 27620 59570 27672 59576
rect 27724 58698 27752 60658
rect 27804 60172 27856 60178
rect 27804 60114 27856 60120
rect 27632 58670 27752 58698
rect 26424 58540 26476 58546
rect 26424 58482 26476 58488
rect 26332 58336 26384 58342
rect 26332 58278 26384 58284
rect 26344 58002 26372 58278
rect 26332 57996 26384 58002
rect 26332 57938 26384 57944
rect 26240 57316 26292 57322
rect 26240 57258 26292 57264
rect 26148 56840 26200 56846
rect 26148 56782 26200 56788
rect 26160 56506 26188 56782
rect 26148 56500 26200 56506
rect 26148 56442 26200 56448
rect 26436 56370 26464 58482
rect 26976 58336 27028 58342
rect 26976 58278 27028 58284
rect 26988 57934 27016 58278
rect 26976 57928 27028 57934
rect 26976 57870 27028 57876
rect 27632 57458 27660 58670
rect 27816 58614 27844 60114
rect 27804 58608 27856 58614
rect 27804 58550 27856 58556
rect 27908 58546 27936 61134
rect 28080 60580 28132 60586
rect 28080 60522 28132 60528
rect 28092 60110 28120 60522
rect 28264 60308 28316 60314
rect 28264 60250 28316 60256
rect 28276 60178 28304 60250
rect 28264 60172 28316 60178
rect 28264 60114 28316 60120
rect 28080 60104 28132 60110
rect 28080 60046 28132 60052
rect 28092 59770 28120 60046
rect 28080 59764 28132 59770
rect 28080 59706 28132 59712
rect 27712 58540 27764 58546
rect 27712 58482 27764 58488
rect 27896 58540 27948 58546
rect 27896 58482 27948 58488
rect 27724 57526 27752 58482
rect 28080 58132 28132 58138
rect 28080 58074 28132 58080
rect 27712 57520 27764 57526
rect 27712 57462 27764 57468
rect 27620 57452 27672 57458
rect 27620 57394 27672 57400
rect 26516 56772 26568 56778
rect 26516 56714 26568 56720
rect 26424 56364 26476 56370
rect 26424 56306 26476 56312
rect 26332 54188 26384 54194
rect 26436 54176 26464 56306
rect 26528 55962 26556 56714
rect 27528 56704 27580 56710
rect 27528 56646 27580 56652
rect 27540 56438 27568 56646
rect 26884 56432 26936 56438
rect 26884 56374 26936 56380
rect 27528 56432 27580 56438
rect 27528 56374 27580 56380
rect 26896 55962 26924 56374
rect 27160 56296 27212 56302
rect 27160 56238 27212 56244
rect 26516 55956 26568 55962
rect 26516 55898 26568 55904
rect 26884 55956 26936 55962
rect 26884 55898 26936 55904
rect 27172 55418 27200 56238
rect 27540 55690 27568 56374
rect 27632 55758 27660 57394
rect 28092 57390 28120 58074
rect 28080 57384 28132 57390
rect 28080 57326 28132 57332
rect 28368 55758 28396 61134
rect 29104 60734 29132 62766
rect 29380 62354 29408 71318
rect 30258 71200 30370 72000
rect 31546 71200 31658 72000
rect 32834 71200 32946 72000
rect 34122 71200 34234 72000
rect 35410 71346 35522 72000
rect 35410 71318 35664 71346
rect 35410 71200 35522 71318
rect 30300 68134 30328 71200
rect 31208 69216 31260 69222
rect 31208 69158 31260 69164
rect 31220 68882 31248 69158
rect 31588 68882 31616 71200
rect 35636 69494 35664 71318
rect 36698 71200 36810 72000
rect 37986 71200 38098 72000
rect 39274 71200 39386 72000
rect 40562 71200 40674 72000
rect 41850 71200 41962 72000
rect 43138 71200 43250 72000
rect 44426 71200 44538 72000
rect 45714 71200 45826 72000
rect 47002 71200 47114 72000
rect 47646 71346 47758 72000
rect 47412 71318 47758 71346
rect 35624 69488 35676 69494
rect 35624 69430 35676 69436
rect 36636 69216 36688 69222
rect 36636 69158 36688 69164
rect 34934 69116 35242 69136
rect 34934 69114 34940 69116
rect 34996 69114 35020 69116
rect 35076 69114 35100 69116
rect 35156 69114 35180 69116
rect 35236 69114 35242 69116
rect 34996 69062 34998 69114
rect 35178 69062 35180 69114
rect 34934 69060 34940 69062
rect 34996 69060 35020 69062
rect 35076 69060 35100 69062
rect 35156 69060 35180 69062
rect 35236 69060 35242 69062
rect 34934 69040 35242 69060
rect 36648 68882 36676 69158
rect 36740 68882 36768 71200
rect 36912 69284 36964 69290
rect 36912 69226 36964 69232
rect 31208 68876 31260 68882
rect 31208 68818 31260 68824
rect 31576 68876 31628 68882
rect 31576 68818 31628 68824
rect 36636 68876 36688 68882
rect 36636 68818 36688 68824
rect 36728 68876 36780 68882
rect 36728 68818 36780 68824
rect 31208 68740 31260 68746
rect 31208 68682 31260 68688
rect 36544 68740 36596 68746
rect 36544 68682 36596 68688
rect 31220 68474 31248 68682
rect 36556 68474 36584 68682
rect 31208 68468 31260 68474
rect 31208 68410 31260 68416
rect 36544 68468 36596 68474
rect 36544 68410 36596 68416
rect 31024 68332 31076 68338
rect 31024 68274 31076 68280
rect 36452 68332 36504 68338
rect 36452 68274 36504 68280
rect 30288 68128 30340 68134
rect 30288 68070 30340 68076
rect 31036 67794 31064 68274
rect 34934 68028 35242 68048
rect 34934 68026 34940 68028
rect 34996 68026 35020 68028
rect 35076 68026 35100 68028
rect 35156 68026 35180 68028
rect 35236 68026 35242 68028
rect 34996 67974 34998 68026
rect 35178 67974 35180 68026
rect 34934 67972 34940 67974
rect 34996 67972 35020 67974
rect 35076 67972 35100 67974
rect 35156 67972 35180 67974
rect 35236 67972 35242 67974
rect 34934 67952 35242 67972
rect 31024 67788 31076 67794
rect 31024 67730 31076 67736
rect 31036 62490 31064 67730
rect 36464 67114 36492 68274
rect 36452 67108 36504 67114
rect 36452 67050 36504 67056
rect 34934 66940 35242 66960
rect 34934 66938 34940 66940
rect 34996 66938 35020 66940
rect 35076 66938 35100 66940
rect 35156 66938 35180 66940
rect 35236 66938 35242 66940
rect 34996 66886 34998 66938
rect 35178 66886 35180 66938
rect 34934 66884 34940 66886
rect 34996 66884 35020 66886
rect 35076 66884 35100 66886
rect 35156 66884 35180 66886
rect 35236 66884 35242 66886
rect 34934 66864 35242 66884
rect 36084 66156 36136 66162
rect 36084 66098 36136 66104
rect 35900 65952 35952 65958
rect 35900 65894 35952 65900
rect 34934 65852 35242 65872
rect 34934 65850 34940 65852
rect 34996 65850 35020 65852
rect 35076 65850 35100 65852
rect 35156 65850 35180 65852
rect 35236 65850 35242 65852
rect 34996 65798 34998 65850
rect 35178 65798 35180 65850
rect 34934 65796 34940 65798
rect 34996 65796 35020 65798
rect 35076 65796 35100 65798
rect 35156 65796 35180 65798
rect 35236 65796 35242 65798
rect 34934 65776 35242 65796
rect 35912 65550 35940 65894
rect 33968 65544 34020 65550
rect 33968 65486 34020 65492
rect 35900 65544 35952 65550
rect 35900 65486 35952 65492
rect 33980 63918 34008 65486
rect 36096 65074 36124 66098
rect 36360 66088 36412 66094
rect 36280 66036 36360 66042
rect 36280 66030 36412 66036
rect 36280 66014 36400 66030
rect 36280 65414 36308 66014
rect 36360 65952 36412 65958
rect 36360 65894 36412 65900
rect 36268 65408 36320 65414
rect 36268 65350 36320 65356
rect 36280 65074 36308 65350
rect 36372 65074 36400 65894
rect 36084 65068 36136 65074
rect 36084 65010 36136 65016
rect 36268 65068 36320 65074
rect 36268 65010 36320 65016
rect 36360 65068 36412 65074
rect 36360 65010 36412 65016
rect 34934 64764 35242 64784
rect 34934 64762 34940 64764
rect 34996 64762 35020 64764
rect 35076 64762 35100 64764
rect 35156 64762 35180 64764
rect 35236 64762 35242 64764
rect 34996 64710 34998 64762
rect 35178 64710 35180 64762
rect 34934 64708 34940 64710
rect 34996 64708 35020 64710
rect 35076 64708 35100 64710
rect 35156 64708 35180 64710
rect 35236 64708 35242 64710
rect 34934 64688 35242 64708
rect 34704 63980 34756 63986
rect 34704 63922 34756 63928
rect 33416 63912 33468 63918
rect 33416 63854 33468 63860
rect 33968 63912 34020 63918
rect 33968 63854 34020 63860
rect 31944 63232 31996 63238
rect 31944 63174 31996 63180
rect 31024 62484 31076 62490
rect 31024 62426 31076 62432
rect 29368 62348 29420 62354
rect 29368 62290 29420 62296
rect 29736 62280 29788 62286
rect 29736 62222 29788 62228
rect 30380 62280 30432 62286
rect 30380 62222 30432 62228
rect 29748 62150 29776 62222
rect 29736 62144 29788 62150
rect 29736 62086 29788 62092
rect 29748 61334 29776 62086
rect 30288 61804 30340 61810
rect 30288 61746 30340 61752
rect 29736 61328 29788 61334
rect 29736 61270 29788 61276
rect 30300 60858 30328 61746
rect 30392 61606 30420 62222
rect 31760 61872 31812 61878
rect 31760 61814 31812 61820
rect 30380 61600 30432 61606
rect 30380 61542 30432 61548
rect 30288 60852 30340 60858
rect 30288 60794 30340 60800
rect 29104 60706 29224 60734
rect 30392 60722 30420 61542
rect 31484 61260 31536 61266
rect 31484 61202 31536 61208
rect 31024 61192 31076 61198
rect 31024 61134 31076 61140
rect 31208 61192 31260 61198
rect 31208 61134 31260 61140
rect 28540 60172 28592 60178
rect 28540 60114 28592 60120
rect 28552 59634 28580 60114
rect 28540 59628 28592 59634
rect 28540 59570 28592 59576
rect 28908 59628 28960 59634
rect 28908 59570 28960 59576
rect 28920 58834 28948 59570
rect 28736 58806 29132 58834
rect 28540 58472 28592 58478
rect 28540 58414 28592 58420
rect 28552 56506 28580 58414
rect 28736 57050 28764 58806
rect 28908 58676 28960 58682
rect 28908 58618 28960 58624
rect 28920 58546 28948 58618
rect 29104 58546 29132 58806
rect 28908 58540 28960 58546
rect 28908 58482 28960 58488
rect 29092 58540 29144 58546
rect 29092 58482 29144 58488
rect 28816 58472 28868 58478
rect 28816 58414 28868 58420
rect 28828 58138 28856 58414
rect 28816 58132 28868 58138
rect 28816 58074 28868 58080
rect 28724 57044 28776 57050
rect 28724 56986 28776 56992
rect 28632 56772 28684 56778
rect 28632 56714 28684 56720
rect 28540 56500 28592 56506
rect 28540 56442 28592 56448
rect 28540 56364 28592 56370
rect 28540 56306 28592 56312
rect 28448 56228 28500 56234
rect 28448 56170 28500 56176
rect 28460 55826 28488 56170
rect 28448 55820 28500 55826
rect 28448 55762 28500 55768
rect 27620 55752 27672 55758
rect 27620 55694 27672 55700
rect 28356 55752 28408 55758
rect 28356 55694 28408 55700
rect 27528 55684 27580 55690
rect 27528 55626 27580 55632
rect 27160 55412 27212 55418
rect 27160 55354 27212 55360
rect 27632 55026 27660 55694
rect 27632 54998 27844 55026
rect 26384 54148 26464 54176
rect 27068 54188 27120 54194
rect 26332 54130 26384 54136
rect 27068 54130 27120 54136
rect 26240 53712 26292 53718
rect 26240 53654 26292 53660
rect 26252 53174 26280 53654
rect 26240 53168 26292 53174
rect 26240 53110 26292 53116
rect 26344 53038 26372 54130
rect 27080 53786 27108 54130
rect 27068 53780 27120 53786
rect 27068 53722 27120 53728
rect 27252 53780 27304 53786
rect 27252 53722 27304 53728
rect 27264 53514 27292 53722
rect 27816 53582 27844 54998
rect 28368 54074 28396 55694
rect 28552 55418 28580 56306
rect 28540 55412 28592 55418
rect 28540 55354 28592 55360
rect 28276 54046 28396 54074
rect 27804 53576 27856 53582
rect 27804 53518 27856 53524
rect 27252 53508 27304 53514
rect 27252 53450 27304 53456
rect 26332 53032 26384 53038
rect 26332 52974 26384 52980
rect 27436 52896 27488 52902
rect 27436 52838 27488 52844
rect 27448 52494 27476 52838
rect 26792 52488 26844 52494
rect 26792 52430 26844 52436
rect 27436 52488 27488 52494
rect 27436 52430 27488 52436
rect 26804 51610 26832 52430
rect 27816 51950 27844 53518
rect 28172 53032 28224 53038
rect 28172 52974 28224 52980
rect 28184 52698 28212 52974
rect 28172 52692 28224 52698
rect 28172 52634 28224 52640
rect 28276 52358 28304 54046
rect 28356 53984 28408 53990
rect 28356 53926 28408 53932
rect 28368 53514 28396 53926
rect 28356 53508 28408 53514
rect 28356 53450 28408 53456
rect 28368 53038 28396 53450
rect 28448 53100 28500 53106
rect 28448 53042 28500 53048
rect 28356 53032 28408 53038
rect 28356 52974 28408 52980
rect 28460 52698 28488 53042
rect 28448 52692 28500 52698
rect 28448 52634 28500 52640
rect 28264 52352 28316 52358
rect 28264 52294 28316 52300
rect 28276 52018 28304 52294
rect 28080 52012 28132 52018
rect 28080 51954 28132 51960
rect 28264 52012 28316 52018
rect 28264 51954 28316 51960
rect 27804 51944 27856 51950
rect 27804 51886 27856 51892
rect 27804 51808 27856 51814
rect 27804 51750 27856 51756
rect 26792 51604 26844 51610
rect 26792 51546 26844 51552
rect 26332 51536 26384 51542
rect 26332 51478 26384 51484
rect 26240 51400 26292 51406
rect 26240 51342 26292 51348
rect 26068 51046 26188 51074
rect 26056 49632 26108 49638
rect 26056 49574 26108 49580
rect 26068 49230 26096 49574
rect 26056 49224 26108 49230
rect 26056 49166 26108 49172
rect 26056 46504 26108 46510
rect 26054 46472 26056 46481
rect 26108 46472 26110 46481
rect 26054 46407 26110 46416
rect 26068 46170 26096 46407
rect 26056 46164 26108 46170
rect 26056 46106 26108 46112
rect 25976 45526 26096 45554
rect 25964 45280 26016 45286
rect 25964 45222 26016 45228
rect 25976 44878 26004 45222
rect 25964 44872 26016 44878
rect 25964 44814 26016 44820
rect 26068 42770 26096 45526
rect 26056 42764 26108 42770
rect 26056 42706 26108 42712
rect 26160 42378 26188 51046
rect 26252 50930 26280 51342
rect 26344 50998 26372 51478
rect 26332 50992 26384 50998
rect 26332 50934 26384 50940
rect 26240 50924 26292 50930
rect 26240 50866 26292 50872
rect 27620 50924 27672 50930
rect 27620 50866 27672 50872
rect 26252 47666 26280 50866
rect 27632 50522 27660 50866
rect 27620 50516 27672 50522
rect 27620 50458 27672 50464
rect 27816 50318 27844 51750
rect 28092 51474 28120 51954
rect 28080 51468 28132 51474
rect 28080 51410 28132 51416
rect 27988 51400 28040 51406
rect 27988 51342 28040 51348
rect 28000 50386 28028 51342
rect 28092 51066 28120 51410
rect 28276 51406 28304 51954
rect 28264 51400 28316 51406
rect 28264 51342 28316 51348
rect 28644 51074 28672 56714
rect 28724 55616 28776 55622
rect 28724 55558 28776 55564
rect 28736 55282 28764 55558
rect 28724 55276 28776 55282
rect 28724 55218 28776 55224
rect 29000 54664 29052 54670
rect 29000 54606 29052 54612
rect 29012 54262 29040 54606
rect 29000 54256 29052 54262
rect 29000 54198 29052 54204
rect 29196 54058 29224 60706
rect 30380 60716 30432 60722
rect 30380 60658 30432 60664
rect 30472 60648 30524 60654
rect 30472 60590 30524 60596
rect 30484 60314 30512 60590
rect 31036 60314 31064 61134
rect 31220 60722 31248 61134
rect 31496 60790 31524 61202
rect 31772 61198 31800 61814
rect 31760 61192 31812 61198
rect 31760 61134 31812 61140
rect 31484 60784 31536 60790
rect 31484 60726 31536 60732
rect 31208 60716 31260 60722
rect 31208 60658 31260 60664
rect 30472 60308 30524 60314
rect 30472 60250 30524 60256
rect 31024 60308 31076 60314
rect 31024 60250 31076 60256
rect 29920 60104 29972 60110
rect 29920 60046 29972 60052
rect 29276 59968 29328 59974
rect 29276 59910 29328 59916
rect 29644 59968 29696 59974
rect 29644 59910 29696 59916
rect 29288 59430 29316 59910
rect 29656 59634 29684 59910
rect 29644 59628 29696 59634
rect 29644 59570 29696 59576
rect 29368 59560 29420 59566
rect 29368 59502 29420 59508
rect 29276 59424 29328 59430
rect 29276 59366 29328 59372
rect 29288 58954 29316 59366
rect 29276 58948 29328 58954
rect 29276 58890 29328 58896
rect 29380 57866 29408 59502
rect 29932 59226 29960 60046
rect 31496 59548 31524 60726
rect 31668 60104 31720 60110
rect 31668 60046 31720 60052
rect 31760 60104 31812 60110
rect 31760 60046 31812 60052
rect 31576 59560 31628 59566
rect 31496 59520 31576 59548
rect 31576 59502 31628 59508
rect 29920 59220 29972 59226
rect 29920 59162 29972 59168
rect 30932 58948 30984 58954
rect 30932 58890 30984 58896
rect 30472 58880 30524 58886
rect 30472 58822 30524 58828
rect 29828 58540 29880 58546
rect 29828 58482 29880 58488
rect 29840 57934 29868 58482
rect 29920 58336 29972 58342
rect 29920 58278 29972 58284
rect 30380 58336 30432 58342
rect 30380 58278 30432 58284
rect 29828 57928 29880 57934
rect 29828 57870 29880 57876
rect 29368 57860 29420 57866
rect 29368 57802 29420 57808
rect 29644 56500 29696 56506
rect 29644 56442 29696 56448
rect 29656 56234 29684 56442
rect 29644 56228 29696 56234
rect 29644 56170 29696 56176
rect 29184 54052 29236 54058
rect 29184 53994 29236 54000
rect 29092 53712 29144 53718
rect 29092 53654 29144 53660
rect 29104 53106 29132 53654
rect 29092 53100 29144 53106
rect 29092 53042 29144 53048
rect 28828 52970 29040 52986
rect 28816 52964 29040 52970
rect 28868 52958 29040 52964
rect 28816 52906 28868 52912
rect 29012 52680 29040 52958
rect 29656 52698 29684 56170
rect 29840 55758 29868 57870
rect 29932 57798 29960 58278
rect 30392 57934 30420 58278
rect 30380 57928 30432 57934
rect 30380 57870 30432 57876
rect 29920 57792 29972 57798
rect 29920 57734 29972 57740
rect 29932 57526 29960 57734
rect 30484 57526 30512 58822
rect 29920 57520 29972 57526
rect 29920 57462 29972 57468
rect 30472 57520 30524 57526
rect 30472 57462 30524 57468
rect 30012 57452 30064 57458
rect 30012 57394 30064 57400
rect 30024 55894 30052 57394
rect 30380 57384 30432 57390
rect 30380 57326 30432 57332
rect 30196 57248 30248 57254
rect 30196 57190 30248 57196
rect 30208 56386 30236 57190
rect 30392 56982 30420 57326
rect 30380 56976 30432 56982
rect 30380 56918 30432 56924
rect 30380 56704 30432 56710
rect 30380 56646 30432 56652
rect 30208 56358 30328 56386
rect 30104 56296 30156 56302
rect 30104 56238 30156 56244
rect 30196 56296 30248 56302
rect 30196 56238 30248 56244
rect 30012 55888 30064 55894
rect 30012 55830 30064 55836
rect 29828 55752 29880 55758
rect 29828 55694 29880 55700
rect 29736 55616 29788 55622
rect 29736 55558 29788 55564
rect 29748 53582 29776 55558
rect 30024 54602 30052 55830
rect 30116 55690 30144 56238
rect 30104 55684 30156 55690
rect 30104 55626 30156 55632
rect 30012 54596 30064 54602
rect 30012 54538 30064 54544
rect 29828 54528 29880 54534
rect 29828 54470 29880 54476
rect 29840 54194 29868 54470
rect 29828 54188 29880 54194
rect 29828 54130 29880 54136
rect 29828 53984 29880 53990
rect 30208 53938 30236 56238
rect 30300 55962 30328 56358
rect 30392 56166 30420 56646
rect 30380 56160 30432 56166
rect 30380 56102 30432 56108
rect 30288 55956 30340 55962
rect 30288 55898 30340 55904
rect 29828 53926 29880 53932
rect 29736 53576 29788 53582
rect 29736 53518 29788 53524
rect 29092 52692 29144 52698
rect 29012 52652 29092 52680
rect 29092 52634 29144 52640
rect 29644 52692 29696 52698
rect 29644 52634 29696 52640
rect 28908 52488 28960 52494
rect 28908 52430 28960 52436
rect 29552 52488 29604 52494
rect 29552 52430 29604 52436
rect 28920 52358 28948 52430
rect 28908 52352 28960 52358
rect 28908 52294 28960 52300
rect 29564 52086 29592 52430
rect 29276 52080 29328 52086
rect 29276 52022 29328 52028
rect 29552 52080 29604 52086
rect 29552 52022 29604 52028
rect 28908 51944 28960 51950
rect 28908 51886 28960 51892
rect 28080 51060 28132 51066
rect 28080 51002 28132 51008
rect 28552 51046 28672 51074
rect 27988 50380 28040 50386
rect 27988 50322 28040 50328
rect 27804 50312 27856 50318
rect 27804 50254 27856 50260
rect 27344 49836 27396 49842
rect 27344 49778 27396 49784
rect 26332 49224 26384 49230
rect 26332 49166 26384 49172
rect 26344 48890 26372 49166
rect 27356 48890 27384 49778
rect 27620 49088 27672 49094
rect 27620 49030 27672 49036
rect 26332 48884 26384 48890
rect 26332 48826 26384 48832
rect 27344 48884 27396 48890
rect 27344 48826 27396 48832
rect 26516 48748 26568 48754
rect 26516 48690 26568 48696
rect 26528 48006 26556 48690
rect 27632 48686 27660 49030
rect 28000 48822 28028 50322
rect 27988 48816 28040 48822
rect 27988 48758 28040 48764
rect 27896 48748 27948 48754
rect 27896 48690 27948 48696
rect 27620 48680 27672 48686
rect 27620 48622 27672 48628
rect 27528 48136 27580 48142
rect 27528 48078 27580 48084
rect 27436 48068 27488 48074
rect 27436 48010 27488 48016
rect 26516 48000 26568 48006
rect 26516 47942 26568 47948
rect 27160 48000 27212 48006
rect 27160 47942 27212 47948
rect 26240 47660 26292 47666
rect 26240 47602 26292 47608
rect 25872 42356 25924 42362
rect 25872 42298 25924 42304
rect 26068 42350 26188 42378
rect 25884 42022 25912 42298
rect 25964 42152 26016 42158
rect 25964 42094 26016 42100
rect 26068 42106 26096 42350
rect 26146 42256 26202 42265
rect 26146 42191 26148 42200
rect 26200 42191 26202 42200
rect 26148 42162 26200 42168
rect 25872 42016 25924 42022
rect 25872 41958 25924 41964
rect 25780 41812 25832 41818
rect 25780 41754 25832 41760
rect 25872 40928 25924 40934
rect 25872 40870 25924 40876
rect 25780 39636 25832 39642
rect 25780 39578 25832 39584
rect 25792 37874 25820 39578
rect 25884 39370 25912 40870
rect 25872 39364 25924 39370
rect 25872 39306 25924 39312
rect 25780 37868 25832 37874
rect 25780 37810 25832 37816
rect 25688 36848 25740 36854
rect 25688 36790 25740 36796
rect 25792 36174 25820 37810
rect 25780 36168 25832 36174
rect 25780 36110 25832 36116
rect 25688 35488 25740 35494
rect 25688 35430 25740 35436
rect 25700 35290 25728 35430
rect 25688 35284 25740 35290
rect 25688 35226 25740 35232
rect 25780 33312 25832 33318
rect 25780 33254 25832 33260
rect 25792 32502 25820 33254
rect 25884 32842 25912 39306
rect 25872 32836 25924 32842
rect 25872 32778 25924 32784
rect 25780 32496 25832 32502
rect 25780 32438 25832 32444
rect 25688 29640 25740 29646
rect 25688 29582 25740 29588
rect 25700 28762 25728 29582
rect 25688 28756 25740 28762
rect 25688 28698 25740 28704
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 25976 2582 26004 42094
rect 26068 42078 26188 42106
rect 26056 42016 26108 42022
rect 26056 41958 26108 41964
rect 26068 40934 26096 41958
rect 26056 40928 26108 40934
rect 26056 40870 26108 40876
rect 26160 40712 26188 42078
rect 26068 40684 26188 40712
rect 26068 39522 26096 40684
rect 26252 40610 26280 47602
rect 26424 47456 26476 47462
rect 26424 47398 26476 47404
rect 26436 47122 26464 47398
rect 26424 47116 26476 47122
rect 26424 47058 26476 47064
rect 26330 46472 26386 46481
rect 26330 46407 26332 46416
rect 26384 46407 26386 46416
rect 26332 46378 26384 46384
rect 26528 45554 26556 47942
rect 27172 47054 27200 47942
rect 27448 47666 27476 48010
rect 27540 47802 27568 48078
rect 27528 47796 27580 47802
rect 27528 47738 27580 47744
rect 27804 47728 27856 47734
rect 27804 47670 27856 47676
rect 27436 47660 27488 47666
rect 27436 47602 27488 47608
rect 27160 47048 27212 47054
rect 27160 46990 27212 46996
rect 27448 45554 27476 47602
rect 27816 47258 27844 47670
rect 27804 47252 27856 47258
rect 27804 47194 27856 47200
rect 26436 45526 26556 45554
rect 27356 45526 27476 45554
rect 26332 41812 26384 41818
rect 26332 41754 26384 41760
rect 26344 41614 26372 41754
rect 26332 41608 26384 41614
rect 26332 41550 26384 41556
rect 26160 40582 26280 40610
rect 26160 39642 26188 40582
rect 26240 40520 26292 40526
rect 26240 40462 26292 40468
rect 26252 40186 26280 40462
rect 26240 40180 26292 40186
rect 26240 40122 26292 40128
rect 26332 40044 26384 40050
rect 26332 39986 26384 39992
rect 26344 39642 26372 39986
rect 26148 39636 26200 39642
rect 26148 39578 26200 39584
rect 26332 39636 26384 39642
rect 26332 39578 26384 39584
rect 26068 39494 26188 39522
rect 26056 37868 26108 37874
rect 26056 37810 26108 37816
rect 26068 34610 26096 37810
rect 26160 37806 26188 39494
rect 26240 39092 26292 39098
rect 26240 39034 26292 39040
rect 26252 38962 26280 39034
rect 26240 38956 26292 38962
rect 26240 38898 26292 38904
rect 26148 37800 26200 37806
rect 26148 37742 26200 37748
rect 26252 36718 26280 38898
rect 26436 37874 26464 45526
rect 26976 45484 27028 45490
rect 26976 45426 27028 45432
rect 26988 44946 27016 45426
rect 26976 44940 27028 44946
rect 26976 44882 27028 44888
rect 27252 44192 27304 44198
rect 27252 44134 27304 44140
rect 27160 43784 27212 43790
rect 27160 43726 27212 43732
rect 26976 43648 27028 43654
rect 26976 43590 27028 43596
rect 26988 43314 27016 43590
rect 27172 43450 27200 43726
rect 27160 43444 27212 43450
rect 27160 43386 27212 43392
rect 27264 43382 27292 44134
rect 27252 43376 27304 43382
rect 27252 43318 27304 43324
rect 26976 43308 27028 43314
rect 26976 43250 27028 43256
rect 26976 42696 27028 42702
rect 26976 42638 27028 42644
rect 26988 42226 27016 42638
rect 26976 42220 27028 42226
rect 26976 42162 27028 42168
rect 26516 41812 26568 41818
rect 26516 41754 26568 41760
rect 26424 37868 26476 37874
rect 26424 37810 26476 37816
rect 26240 36712 26292 36718
rect 26240 36654 26292 36660
rect 26056 34604 26108 34610
rect 26056 34546 26108 34552
rect 26068 32434 26096 34546
rect 26240 32904 26292 32910
rect 26240 32846 26292 32852
rect 26252 32570 26280 32846
rect 26240 32564 26292 32570
rect 26240 32506 26292 32512
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 26068 31822 26096 32370
rect 26056 31816 26108 31822
rect 26056 31758 26108 31764
rect 26528 31754 26556 41754
rect 27252 40996 27304 41002
rect 27252 40938 27304 40944
rect 26976 40452 27028 40458
rect 26976 40394 27028 40400
rect 26988 40186 27016 40394
rect 26976 40180 27028 40186
rect 26976 40122 27028 40128
rect 27264 39642 27292 40938
rect 27252 39636 27304 39642
rect 27252 39578 27304 39584
rect 27264 39438 27292 39578
rect 26792 39432 26844 39438
rect 26792 39374 26844 39380
rect 27252 39432 27304 39438
rect 27252 39374 27304 39380
rect 26608 37188 26660 37194
rect 26608 37130 26660 37136
rect 26620 36378 26648 37130
rect 26608 36372 26660 36378
rect 26608 36314 26660 36320
rect 26700 31816 26752 31822
rect 26700 31758 26752 31764
rect 26436 31726 26556 31754
rect 26332 31136 26384 31142
rect 26332 31078 26384 31084
rect 26344 30938 26372 31078
rect 26332 30932 26384 30938
rect 26332 30874 26384 30880
rect 26056 29504 26108 29510
rect 26056 29446 26108 29452
rect 26068 28966 26096 29446
rect 26056 28960 26108 28966
rect 26056 28902 26108 28908
rect 26068 28626 26096 28902
rect 26056 28620 26108 28626
rect 26056 28562 26108 28568
rect 26332 28416 26384 28422
rect 26332 28358 26384 28364
rect 26148 27532 26200 27538
rect 26148 27474 26200 27480
rect 26160 3398 26188 27474
rect 26344 26994 26372 28358
rect 26332 26988 26384 26994
rect 26332 26930 26384 26936
rect 26436 26234 26464 31726
rect 26516 31680 26568 31686
rect 26516 31622 26568 31628
rect 26528 31414 26556 31622
rect 26712 31482 26740 31758
rect 26700 31476 26752 31482
rect 26700 31418 26752 31424
rect 26516 31408 26568 31414
rect 26516 31350 26568 31356
rect 26516 31136 26568 31142
rect 26516 31078 26568 31084
rect 26528 29714 26556 31078
rect 26804 30938 26832 39374
rect 27068 39296 27120 39302
rect 27068 39238 27120 39244
rect 27080 38962 27108 39238
rect 27356 39098 27384 45526
rect 27620 45416 27672 45422
rect 27620 45358 27672 45364
rect 27632 45082 27660 45358
rect 27620 45076 27672 45082
rect 27620 45018 27672 45024
rect 27528 42220 27580 42226
rect 27528 42162 27580 42168
rect 27540 41818 27568 42162
rect 27528 41812 27580 41818
rect 27528 41754 27580 41760
rect 27712 41608 27764 41614
rect 27712 41550 27764 41556
rect 27724 41206 27752 41550
rect 27908 41414 27936 48690
rect 28448 48680 28500 48686
rect 28448 48622 28500 48628
rect 28460 47666 28488 48622
rect 28552 47734 28580 51046
rect 28920 50862 28948 51886
rect 28908 50856 28960 50862
rect 28908 50798 28960 50804
rect 29184 49836 29236 49842
rect 29184 49778 29236 49784
rect 28632 49632 28684 49638
rect 28632 49574 28684 49580
rect 28644 49230 28672 49574
rect 28724 49360 28776 49366
rect 28724 49302 28776 49308
rect 28632 49224 28684 49230
rect 28632 49166 28684 49172
rect 28736 48754 28764 49302
rect 29092 49088 29144 49094
rect 29092 49030 29144 49036
rect 29104 48822 29132 49030
rect 29196 48890 29224 49778
rect 29184 48884 29236 48890
rect 29184 48826 29236 48832
rect 29092 48816 29144 48822
rect 29092 48758 29144 48764
rect 28724 48748 28776 48754
rect 28724 48690 28776 48696
rect 29104 47734 29132 48758
rect 29184 48000 29236 48006
rect 29184 47942 29236 47948
rect 28540 47728 28592 47734
rect 28540 47670 28592 47676
rect 29092 47728 29144 47734
rect 29092 47670 29144 47676
rect 28448 47660 28500 47666
rect 28448 47602 28500 47608
rect 27988 46572 28040 46578
rect 27988 46514 28040 46520
rect 27816 41386 27936 41414
rect 27712 41200 27764 41206
rect 27712 41142 27764 41148
rect 27816 39982 27844 41386
rect 27804 39976 27856 39982
rect 27804 39918 27856 39924
rect 27344 39092 27396 39098
rect 27344 39034 27396 39040
rect 27068 38956 27120 38962
rect 27068 38898 27120 38904
rect 27712 38956 27764 38962
rect 27712 38898 27764 38904
rect 27724 38554 27752 38898
rect 27712 38548 27764 38554
rect 27712 38490 27764 38496
rect 27252 38208 27304 38214
rect 27252 38150 27304 38156
rect 27160 37936 27212 37942
rect 27160 37878 27212 37884
rect 27172 37330 27200 37878
rect 27264 37466 27292 38150
rect 27344 37664 27396 37670
rect 27344 37606 27396 37612
rect 27528 37664 27580 37670
rect 27528 37606 27580 37612
rect 27252 37460 27304 37466
rect 27252 37402 27304 37408
rect 27264 37330 27292 37402
rect 27160 37324 27212 37330
rect 27160 37266 27212 37272
rect 27252 37324 27304 37330
rect 27252 37266 27304 37272
rect 27356 36718 27384 37606
rect 27344 36712 27396 36718
rect 27344 36654 27396 36660
rect 26976 35488 27028 35494
rect 26976 35430 27028 35436
rect 26988 35086 27016 35430
rect 27068 35148 27120 35154
rect 27068 35090 27120 35096
rect 26976 35080 27028 35086
rect 26976 35022 27028 35028
rect 27080 34678 27108 35090
rect 27068 34672 27120 34678
rect 27068 34614 27120 34620
rect 27356 34406 27384 36654
rect 27540 36174 27568 37606
rect 27712 37392 27764 37398
rect 27712 37334 27764 37340
rect 27528 36168 27580 36174
rect 27528 36110 27580 36116
rect 27436 35692 27488 35698
rect 27436 35634 27488 35640
rect 27448 34746 27476 35634
rect 27724 35222 27752 37334
rect 27712 35216 27764 35222
rect 27712 35158 27764 35164
rect 27436 34740 27488 34746
rect 27436 34682 27488 34688
rect 27344 34400 27396 34406
rect 27344 34342 27396 34348
rect 27724 33454 27752 35158
rect 27712 33448 27764 33454
rect 27712 33390 27764 33396
rect 27620 33380 27672 33386
rect 27620 33322 27672 33328
rect 27632 33114 27660 33322
rect 27620 33108 27672 33114
rect 27620 33050 27672 33056
rect 27632 32842 27660 33050
rect 26976 32836 27028 32842
rect 26976 32778 27028 32784
rect 27620 32836 27672 32842
rect 27620 32778 27672 32784
rect 26988 32570 27016 32778
rect 27712 32768 27764 32774
rect 27712 32710 27764 32716
rect 26976 32564 27028 32570
rect 26976 32506 27028 32512
rect 27724 31482 27752 32710
rect 27816 31890 27844 39918
rect 27896 39296 27948 39302
rect 27896 39238 27948 39244
rect 27908 38350 27936 39238
rect 27896 38344 27948 38350
rect 27896 38286 27948 38292
rect 28000 37482 28028 46514
rect 28356 45824 28408 45830
rect 28356 45766 28408 45772
rect 28368 45558 28396 45766
rect 28356 45552 28408 45558
rect 28356 45494 28408 45500
rect 28356 44872 28408 44878
rect 28356 44814 28408 44820
rect 28368 44198 28396 44814
rect 28356 44192 28408 44198
rect 28356 44134 28408 44140
rect 28368 43790 28396 44134
rect 28080 43784 28132 43790
rect 28356 43784 28408 43790
rect 28080 43726 28132 43732
rect 28276 43744 28356 43772
rect 28092 40594 28120 43726
rect 28276 42242 28304 43744
rect 28356 43726 28408 43732
rect 28356 42764 28408 42770
rect 28356 42706 28408 42712
rect 28368 42362 28396 42706
rect 28356 42356 28408 42362
rect 28356 42298 28408 42304
rect 28276 42214 28396 42242
rect 28172 41608 28224 41614
rect 28170 41576 28172 41585
rect 28224 41576 28226 41585
rect 28170 41511 28226 41520
rect 28264 41064 28316 41070
rect 28264 41006 28316 41012
rect 28080 40588 28132 40594
rect 28080 40530 28132 40536
rect 28276 40526 28304 41006
rect 28264 40520 28316 40526
rect 28264 40462 28316 40468
rect 28276 40050 28304 40462
rect 28264 40044 28316 40050
rect 28264 39986 28316 39992
rect 28276 39438 28304 39986
rect 28172 39432 28224 39438
rect 28172 39374 28224 39380
rect 28264 39432 28316 39438
rect 28264 39374 28316 39380
rect 28184 39098 28212 39374
rect 28172 39092 28224 39098
rect 28172 39034 28224 39040
rect 28368 37482 28396 42214
rect 28448 41132 28500 41138
rect 28448 41074 28500 41080
rect 28460 40934 28488 41074
rect 28448 40928 28500 40934
rect 28448 40870 28500 40876
rect 28448 40384 28500 40390
rect 28448 40326 28500 40332
rect 28460 40118 28488 40326
rect 28448 40112 28500 40118
rect 28448 40054 28500 40060
rect 27908 37454 28028 37482
rect 28276 37454 28396 37482
rect 27908 37398 27936 37454
rect 27896 37392 27948 37398
rect 27896 37334 27948 37340
rect 28080 37256 28132 37262
rect 28080 37198 28132 37204
rect 28092 36242 28120 37198
rect 28080 36236 28132 36242
rect 28080 36178 28132 36184
rect 28080 35080 28132 35086
rect 28080 35022 28132 35028
rect 28092 34202 28120 35022
rect 28172 34400 28224 34406
rect 28172 34342 28224 34348
rect 28080 34196 28132 34202
rect 28080 34138 28132 34144
rect 28184 33114 28212 34342
rect 28276 33998 28304 37454
rect 28552 37346 28580 47670
rect 28908 47592 28960 47598
rect 28908 47534 28960 47540
rect 28920 46918 28948 47534
rect 28908 46912 28960 46918
rect 28908 46854 28960 46860
rect 28632 46708 28684 46714
rect 28632 46650 28684 46656
rect 28644 46374 28672 46650
rect 28920 46578 28948 46854
rect 28908 46572 28960 46578
rect 28908 46514 28960 46520
rect 28632 46368 28684 46374
rect 28632 46310 28684 46316
rect 29000 46368 29052 46374
rect 29000 46310 29052 46316
rect 28908 45892 28960 45898
rect 28908 45834 28960 45840
rect 28816 45552 28868 45558
rect 28816 45494 28868 45500
rect 28828 45286 28856 45494
rect 28816 45280 28868 45286
rect 28816 45222 28868 45228
rect 28828 43654 28856 45222
rect 28920 45082 28948 45834
rect 28908 45076 28960 45082
rect 28908 45018 28960 45024
rect 28908 44396 28960 44402
rect 28908 44338 28960 44344
rect 28920 43926 28948 44338
rect 29012 43994 29040 46310
rect 29000 43988 29052 43994
rect 29000 43930 29052 43936
rect 28908 43920 28960 43926
rect 28908 43862 28960 43868
rect 28816 43648 28868 43654
rect 28816 43590 28868 43596
rect 29012 43314 29040 43930
rect 29000 43308 29052 43314
rect 29000 43250 29052 43256
rect 28632 42220 28684 42226
rect 28632 42162 28684 42168
rect 29092 42220 29144 42226
rect 29092 42162 29144 42168
rect 28368 37318 28580 37346
rect 28368 37262 28396 37318
rect 28356 37256 28408 37262
rect 28356 37198 28408 37204
rect 28368 35086 28396 37198
rect 28448 36168 28500 36174
rect 28448 36110 28500 36116
rect 28356 35080 28408 35086
rect 28356 35022 28408 35028
rect 28368 34202 28396 35022
rect 28356 34196 28408 34202
rect 28356 34138 28408 34144
rect 28264 33992 28316 33998
rect 28264 33934 28316 33940
rect 28264 33448 28316 33454
rect 28264 33390 28316 33396
rect 28356 33448 28408 33454
rect 28356 33390 28408 33396
rect 28460 33402 28488 36110
rect 28540 34196 28592 34202
rect 28540 34138 28592 34144
rect 28552 33522 28580 34138
rect 28540 33516 28592 33522
rect 28540 33458 28592 33464
rect 28172 33108 28224 33114
rect 28172 33050 28224 33056
rect 27804 31884 27856 31890
rect 27804 31826 27856 31832
rect 27712 31476 27764 31482
rect 27712 31418 27764 31424
rect 27804 31408 27856 31414
rect 27804 31350 27856 31356
rect 26792 30932 26844 30938
rect 26792 30874 26844 30880
rect 27816 30054 27844 31350
rect 28080 31136 28132 31142
rect 28184 31124 28212 33050
rect 28276 32298 28304 33390
rect 28368 33318 28396 33390
rect 28460 33374 28580 33402
rect 28356 33312 28408 33318
rect 28356 33254 28408 33260
rect 28448 32768 28500 32774
rect 28448 32710 28500 32716
rect 28460 32434 28488 32710
rect 28448 32428 28500 32434
rect 28448 32370 28500 32376
rect 28264 32292 28316 32298
rect 28264 32234 28316 32240
rect 28552 31822 28580 33374
rect 28540 31816 28592 31822
rect 28540 31758 28592 31764
rect 28132 31096 28212 31124
rect 28540 31136 28592 31142
rect 28080 31078 28132 31084
rect 28540 31078 28592 31084
rect 28552 30734 28580 31078
rect 28540 30728 28592 30734
rect 28540 30670 28592 30676
rect 28356 30592 28408 30598
rect 28356 30534 28408 30540
rect 28368 30326 28396 30534
rect 28356 30320 28408 30326
rect 28356 30262 28408 30268
rect 28080 30116 28132 30122
rect 28080 30058 28132 30064
rect 27344 30048 27396 30054
rect 27344 29990 27396 29996
rect 27804 30048 27856 30054
rect 27804 29990 27856 29996
rect 26516 29708 26568 29714
rect 26516 29650 26568 29656
rect 27356 29646 27384 29990
rect 27712 29844 27764 29850
rect 27712 29786 27764 29792
rect 27344 29640 27396 29646
rect 27344 29582 27396 29588
rect 27620 29504 27672 29510
rect 27620 29446 27672 29452
rect 27436 29096 27488 29102
rect 27436 29038 27488 29044
rect 27448 28014 27476 29038
rect 27632 28150 27660 29446
rect 27724 29016 27752 29786
rect 27816 29306 27844 29990
rect 27804 29300 27856 29306
rect 27804 29242 27856 29248
rect 27896 29300 27948 29306
rect 27896 29242 27948 29248
rect 27804 29028 27856 29034
rect 27724 28988 27804 29016
rect 27908 29016 27936 29242
rect 28092 29170 28120 30058
rect 28080 29164 28132 29170
rect 28080 29106 28132 29112
rect 27856 28988 27936 29016
rect 27804 28970 27856 28976
rect 27620 28144 27672 28150
rect 27620 28086 27672 28092
rect 26516 28008 26568 28014
rect 26516 27950 26568 27956
rect 27436 28008 27488 28014
rect 27436 27950 27488 27956
rect 26528 27130 26556 27950
rect 26608 27872 26660 27878
rect 26608 27814 26660 27820
rect 26516 27124 26568 27130
rect 26516 27066 26568 27072
rect 26620 27062 26648 27814
rect 27632 27674 27660 28086
rect 28356 27872 28408 27878
rect 28356 27814 28408 27820
rect 27620 27668 27672 27674
rect 27620 27610 27672 27616
rect 26976 27464 27028 27470
rect 26976 27406 27028 27412
rect 26988 27130 27016 27406
rect 27528 27396 27580 27402
rect 27528 27338 27580 27344
rect 27620 27396 27672 27402
rect 27620 27338 27672 27344
rect 26976 27124 27028 27130
rect 26976 27066 27028 27072
rect 26608 27056 26660 27062
rect 26608 26998 26660 27004
rect 27540 26586 27568 27338
rect 27632 26994 27660 27338
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 27528 26580 27580 26586
rect 27528 26522 27580 26528
rect 28368 26382 28396 27814
rect 28356 26376 28408 26382
rect 28356 26318 28408 26324
rect 28644 26234 28672 42162
rect 28908 42016 28960 42022
rect 28908 41958 28960 41964
rect 28920 41546 28948 41958
rect 29000 41744 29052 41750
rect 29000 41686 29052 41692
rect 28908 41540 28960 41546
rect 28908 41482 28960 41488
rect 29012 40934 29040 41686
rect 29104 41274 29132 42162
rect 29196 42158 29224 47942
rect 29288 47274 29316 52022
rect 29368 51944 29420 51950
rect 29368 51886 29420 51892
rect 29380 48278 29408 51886
rect 29656 51474 29684 52634
rect 29748 52018 29776 53518
rect 29840 53514 29868 53926
rect 29932 53910 30236 53938
rect 29828 53508 29880 53514
rect 29828 53450 29880 53456
rect 29840 52902 29868 53450
rect 29932 53038 29960 53910
rect 30300 53786 30328 55898
rect 30392 55690 30420 56102
rect 30380 55684 30432 55690
rect 30380 55626 30432 55632
rect 30484 55622 30512 57462
rect 30840 56840 30892 56846
rect 30840 56782 30892 56788
rect 30852 55962 30880 56782
rect 30944 56506 30972 58890
rect 31300 58540 31352 58546
rect 31300 58482 31352 58488
rect 31116 58336 31168 58342
rect 31116 58278 31168 58284
rect 31128 57934 31156 58278
rect 31116 57928 31168 57934
rect 31116 57870 31168 57876
rect 31312 57322 31340 58482
rect 31588 57390 31616 59502
rect 31680 59022 31708 60046
rect 31772 59702 31800 60046
rect 31852 59968 31904 59974
rect 31852 59910 31904 59916
rect 31760 59696 31812 59702
rect 31760 59638 31812 59644
rect 31864 59548 31892 59910
rect 31772 59520 31892 59548
rect 31668 59016 31720 59022
rect 31668 58958 31720 58964
rect 31680 58546 31708 58958
rect 31772 58886 31800 59520
rect 31760 58880 31812 58886
rect 31760 58822 31812 58828
rect 31772 58682 31800 58822
rect 31760 58676 31812 58682
rect 31760 58618 31812 58624
rect 31668 58540 31720 58546
rect 31668 58482 31720 58488
rect 31576 57384 31628 57390
rect 31576 57326 31628 57332
rect 31300 57316 31352 57322
rect 31300 57258 31352 57264
rect 31392 56772 31444 56778
rect 31392 56714 31444 56720
rect 30932 56500 30984 56506
rect 30932 56442 30984 56448
rect 30840 55956 30892 55962
rect 30840 55898 30892 55904
rect 30564 55752 30616 55758
rect 30564 55694 30616 55700
rect 30472 55616 30524 55622
rect 30472 55558 30524 55564
rect 30576 54670 30604 55694
rect 30748 55616 30800 55622
rect 30748 55558 30800 55564
rect 30760 55282 30788 55558
rect 31404 55418 31432 56714
rect 31392 55412 31444 55418
rect 31392 55354 31444 55360
rect 30748 55276 30800 55282
rect 30748 55218 30800 55224
rect 31680 54738 31708 58482
rect 31668 54732 31720 54738
rect 31668 54674 31720 54680
rect 31772 54670 31800 58618
rect 30564 54664 30616 54670
rect 30564 54606 30616 54612
rect 31760 54664 31812 54670
rect 31760 54606 31812 54612
rect 31852 54664 31904 54670
rect 31852 54606 31904 54612
rect 30012 53780 30064 53786
rect 30012 53722 30064 53728
rect 30288 53780 30340 53786
rect 30288 53722 30340 53728
rect 29920 53032 29972 53038
rect 29920 52974 29972 52980
rect 29828 52896 29880 52902
rect 29828 52838 29880 52844
rect 29736 52012 29788 52018
rect 29736 51954 29788 51960
rect 30024 51814 30052 53722
rect 30104 53712 30156 53718
rect 30104 53654 30156 53660
rect 30116 53446 30144 53654
rect 30104 53440 30156 53446
rect 30104 53382 30156 53388
rect 30576 52630 30604 54606
rect 30656 54188 30708 54194
rect 30656 54130 30708 54136
rect 30668 53786 30696 54130
rect 30656 53780 30708 53786
rect 30656 53722 30708 53728
rect 31772 53650 31800 54606
rect 31760 53644 31812 53650
rect 31760 53586 31812 53592
rect 31864 53242 31892 54606
rect 31852 53236 31904 53242
rect 31852 53178 31904 53184
rect 30748 53032 30800 53038
rect 30748 52974 30800 52980
rect 30564 52624 30616 52630
rect 30564 52566 30616 52572
rect 30380 52488 30432 52494
rect 30380 52430 30432 52436
rect 30012 51808 30064 51814
rect 30012 51750 30064 51756
rect 29644 51468 29696 51474
rect 29644 51410 29696 51416
rect 29552 50788 29604 50794
rect 29552 50730 29604 50736
rect 29564 48822 29592 50730
rect 29736 50448 29788 50454
rect 29736 50390 29788 50396
rect 29748 49774 29776 50390
rect 30024 50318 30052 51750
rect 29920 50312 29972 50318
rect 29920 50254 29972 50260
rect 30012 50312 30064 50318
rect 30012 50254 30064 50260
rect 30288 50312 30340 50318
rect 30288 50254 30340 50260
rect 29932 50182 29960 50254
rect 29920 50176 29972 50182
rect 29920 50118 29972 50124
rect 29736 49768 29788 49774
rect 29736 49710 29788 49716
rect 29552 48816 29604 48822
rect 29552 48758 29604 48764
rect 29368 48272 29420 48278
rect 29368 48214 29420 48220
rect 29460 47456 29512 47462
rect 29460 47398 29512 47404
rect 29288 47246 29408 47274
rect 29276 47116 29328 47122
rect 29276 47058 29328 47064
rect 29288 46578 29316 47058
rect 29276 46572 29328 46578
rect 29276 46514 29328 46520
rect 29380 46374 29408 47246
rect 29368 46368 29420 46374
rect 29368 46310 29420 46316
rect 29368 45892 29420 45898
rect 29368 45834 29420 45840
rect 29380 45626 29408 45834
rect 29368 45620 29420 45626
rect 29368 45562 29420 45568
rect 29472 43466 29500 47398
rect 29564 43874 29592 48758
rect 29748 44010 29776 49710
rect 30024 48550 30052 50254
rect 30300 49858 30328 50254
rect 30116 49842 30328 49858
rect 30104 49836 30328 49842
rect 30156 49830 30328 49836
rect 30104 49778 30156 49784
rect 30300 49230 30328 49830
rect 30288 49224 30340 49230
rect 30288 49166 30340 49172
rect 30300 48822 30328 49166
rect 30288 48816 30340 48822
rect 30288 48758 30340 48764
rect 30104 48612 30156 48618
rect 30104 48554 30156 48560
rect 30012 48544 30064 48550
rect 30012 48486 30064 48492
rect 30012 46572 30064 46578
rect 30012 46514 30064 46520
rect 29920 46368 29972 46374
rect 29920 46310 29972 46316
rect 29932 46034 29960 46310
rect 29920 46028 29972 46034
rect 29920 45970 29972 45976
rect 29828 45960 29880 45966
rect 29828 45902 29880 45908
rect 29840 45626 29868 45902
rect 29828 45620 29880 45626
rect 29828 45562 29880 45568
rect 30024 44946 30052 46514
rect 30012 44940 30064 44946
rect 30012 44882 30064 44888
rect 30012 44804 30064 44810
rect 30012 44746 30064 44752
rect 29920 44532 29972 44538
rect 29920 44474 29972 44480
rect 29748 43982 29868 44010
rect 29564 43846 29776 43874
rect 29552 43716 29604 43722
rect 29552 43658 29604 43664
rect 29288 43438 29500 43466
rect 29564 43450 29592 43658
rect 29552 43444 29604 43450
rect 29184 42152 29236 42158
rect 29184 42094 29236 42100
rect 29184 42016 29236 42022
rect 29184 41958 29236 41964
rect 29196 41478 29224 41958
rect 29184 41472 29236 41478
rect 29184 41414 29236 41420
rect 29092 41268 29144 41274
rect 29092 41210 29144 41216
rect 29092 41132 29144 41138
rect 29092 41074 29144 41080
rect 29104 41002 29132 41074
rect 29092 40996 29144 41002
rect 29092 40938 29144 40944
rect 29000 40928 29052 40934
rect 29000 40870 29052 40876
rect 29104 40526 29132 40938
rect 29288 40594 29316 43438
rect 29552 43386 29604 43392
rect 29644 43444 29696 43450
rect 29644 43386 29696 43392
rect 29656 43330 29684 43386
rect 29564 43314 29684 43330
rect 29552 43308 29684 43314
rect 29604 43302 29684 43308
rect 29552 43250 29604 43256
rect 29460 43240 29512 43246
rect 29748 43194 29776 43846
rect 29460 43182 29512 43188
rect 29368 42152 29420 42158
rect 29368 42094 29420 42100
rect 29276 40588 29328 40594
rect 29276 40530 29328 40536
rect 29092 40520 29144 40526
rect 29092 40462 29144 40468
rect 29276 40384 29328 40390
rect 29276 40326 29328 40332
rect 29288 40050 29316 40326
rect 29276 40044 29328 40050
rect 29276 39986 29328 39992
rect 28816 37936 28868 37942
rect 28816 37878 28868 37884
rect 28828 36718 28856 37878
rect 29380 37874 29408 42094
rect 29472 41750 29500 43182
rect 29564 43166 29776 43194
rect 29564 42702 29592 43166
rect 29552 42696 29604 42702
rect 29552 42638 29604 42644
rect 29460 41744 29512 41750
rect 29460 41686 29512 41692
rect 29368 37868 29420 37874
rect 29368 37810 29420 37816
rect 28816 36712 28868 36718
rect 28816 36654 28868 36660
rect 28724 36032 28776 36038
rect 28724 35974 28776 35980
rect 28736 35698 28764 35974
rect 28724 35692 28776 35698
rect 28724 35634 28776 35640
rect 28828 34678 28856 36654
rect 29564 36650 29592 42638
rect 29736 42628 29788 42634
rect 29736 42570 29788 42576
rect 29748 42362 29776 42570
rect 29736 42356 29788 42362
rect 29736 42298 29788 42304
rect 29840 39574 29868 43982
rect 29932 43722 29960 44474
rect 29920 43716 29972 43722
rect 29920 43658 29972 43664
rect 29932 42634 29960 43658
rect 29920 42628 29972 42634
rect 29920 42570 29972 42576
rect 29920 41608 29972 41614
rect 29920 41550 29972 41556
rect 29932 41274 29960 41550
rect 29920 41268 29972 41274
rect 29920 41210 29972 41216
rect 29828 39568 29880 39574
rect 29828 39510 29880 39516
rect 29644 38208 29696 38214
rect 29644 38150 29696 38156
rect 29656 37942 29684 38150
rect 29644 37936 29696 37942
rect 29644 37878 29696 37884
rect 30024 37670 30052 44746
rect 30116 42090 30144 48554
rect 30392 48278 30420 52430
rect 30472 51400 30524 51406
rect 30472 51342 30524 51348
rect 30484 51066 30512 51342
rect 30472 51060 30524 51066
rect 30472 51002 30524 51008
rect 30576 50930 30604 52566
rect 30760 51474 30788 52974
rect 31392 52964 31444 52970
rect 31392 52906 31444 52912
rect 31208 52896 31260 52902
rect 31208 52838 31260 52844
rect 31220 52494 31248 52838
rect 31404 52698 31432 52906
rect 31392 52692 31444 52698
rect 31392 52634 31444 52640
rect 31116 52488 31168 52494
rect 31116 52430 31168 52436
rect 31208 52488 31260 52494
rect 31208 52430 31260 52436
rect 30748 51468 30800 51474
rect 30748 51410 30800 51416
rect 30760 51074 30788 51410
rect 30668 51046 30788 51074
rect 30564 50924 30616 50930
rect 30564 50866 30616 50872
rect 30288 48272 30340 48278
rect 30288 48214 30340 48220
rect 30380 48272 30432 48278
rect 30380 48214 30432 48220
rect 30300 48113 30328 48214
rect 30564 48136 30616 48142
rect 30286 48104 30342 48113
rect 30564 48078 30616 48084
rect 30286 48039 30342 48048
rect 30196 48000 30248 48006
rect 30196 47942 30248 47948
rect 30208 47666 30236 47942
rect 30196 47660 30248 47666
rect 30196 47602 30248 47608
rect 30196 47456 30248 47462
rect 30196 47398 30248 47404
rect 30208 46986 30236 47398
rect 30576 47258 30604 48078
rect 30380 47252 30432 47258
rect 30380 47194 30432 47200
rect 30564 47252 30616 47258
rect 30564 47194 30616 47200
rect 30288 47184 30340 47190
rect 30288 47126 30340 47132
rect 30300 46986 30328 47126
rect 30392 47002 30420 47194
rect 30392 46986 30604 47002
rect 30196 46980 30248 46986
rect 30196 46922 30248 46928
rect 30288 46980 30340 46986
rect 30288 46922 30340 46928
rect 30392 46980 30616 46986
rect 30392 46974 30564 46980
rect 30300 44810 30328 46922
rect 30288 44804 30340 44810
rect 30288 44746 30340 44752
rect 30196 43240 30248 43246
rect 30196 43182 30248 43188
rect 30208 42566 30236 43182
rect 30196 42560 30248 42566
rect 30196 42502 30248 42508
rect 30104 42084 30156 42090
rect 30104 42026 30156 42032
rect 30196 38344 30248 38350
rect 30196 38286 30248 38292
rect 30012 37664 30064 37670
rect 30012 37606 30064 37612
rect 30024 37398 30052 37606
rect 30012 37392 30064 37398
rect 30012 37334 30064 37340
rect 30012 37256 30064 37262
rect 30012 37198 30064 37204
rect 29828 37120 29880 37126
rect 29828 37062 29880 37068
rect 29736 36916 29788 36922
rect 29736 36858 29788 36864
rect 29552 36644 29604 36650
rect 29552 36586 29604 36592
rect 29552 36032 29604 36038
rect 29552 35974 29604 35980
rect 29564 35766 29592 35974
rect 29552 35760 29604 35766
rect 29552 35702 29604 35708
rect 29748 34950 29776 36858
rect 29840 36854 29868 37062
rect 30024 36922 30052 37198
rect 30208 36922 30236 38286
rect 30392 37754 30420 46974
rect 30564 46922 30616 46928
rect 30472 45824 30524 45830
rect 30472 45766 30524 45772
rect 30484 45558 30512 45766
rect 30472 45552 30524 45558
rect 30472 45494 30524 45500
rect 30564 45552 30616 45558
rect 30564 45494 30616 45500
rect 30484 43450 30512 45494
rect 30576 45014 30604 45494
rect 30668 45082 30696 51046
rect 31128 50998 31156 52430
rect 31208 51876 31260 51882
rect 31208 51818 31260 51824
rect 31220 50998 31248 51818
rect 31392 51060 31444 51066
rect 31392 51002 31444 51008
rect 31116 50992 31168 50998
rect 31116 50934 31168 50940
rect 31208 50992 31260 50998
rect 31208 50934 31260 50940
rect 31300 50720 31352 50726
rect 31300 50662 31352 50668
rect 30932 49836 30984 49842
rect 30932 49778 30984 49784
rect 30944 49434 30972 49778
rect 30932 49428 30984 49434
rect 30932 49370 30984 49376
rect 31312 49230 31340 50662
rect 31404 49774 31432 51002
rect 31392 49768 31444 49774
rect 31392 49710 31444 49716
rect 31300 49224 31352 49230
rect 31300 49166 31352 49172
rect 30840 49156 30892 49162
rect 30840 49098 30892 49104
rect 30748 46368 30800 46374
rect 30748 46310 30800 46316
rect 30760 45966 30788 46310
rect 30748 45960 30800 45966
rect 30748 45902 30800 45908
rect 30656 45076 30708 45082
rect 30656 45018 30708 45024
rect 30564 45008 30616 45014
rect 30564 44950 30616 44956
rect 30748 44464 30800 44470
rect 30748 44406 30800 44412
rect 30564 44192 30616 44198
rect 30564 44134 30616 44140
rect 30472 43444 30524 43450
rect 30472 43386 30524 43392
rect 30576 43246 30604 44134
rect 30760 43654 30788 44406
rect 30748 43648 30800 43654
rect 30748 43590 30800 43596
rect 30564 43240 30616 43246
rect 30564 43182 30616 43188
rect 30760 43110 30788 43590
rect 30748 43104 30800 43110
rect 30748 43046 30800 43052
rect 30748 42696 30800 42702
rect 30852 42650 30880 49098
rect 31576 48272 31628 48278
rect 31576 48214 31628 48220
rect 31116 48000 31168 48006
rect 31116 47942 31168 47948
rect 31128 47734 31156 47942
rect 31116 47728 31168 47734
rect 31116 47670 31168 47676
rect 31588 47054 31616 48214
rect 31576 47048 31628 47054
rect 31576 46990 31628 46996
rect 31852 46912 31904 46918
rect 31852 46854 31904 46860
rect 30932 46572 30984 46578
rect 30932 46514 30984 46520
rect 30944 45626 30972 46514
rect 31864 46510 31892 46854
rect 31852 46504 31904 46510
rect 31852 46446 31904 46452
rect 30932 45620 30984 45626
rect 30932 45562 30984 45568
rect 31116 44872 31168 44878
rect 31116 44814 31168 44820
rect 30932 44736 30984 44742
rect 30932 44678 30984 44684
rect 30944 43858 30972 44678
rect 30932 43852 30984 43858
rect 30932 43794 30984 43800
rect 31024 43240 31076 43246
rect 31024 43182 31076 43188
rect 31036 42906 31064 43182
rect 31024 42900 31076 42906
rect 31024 42842 31076 42848
rect 30800 42644 30880 42650
rect 30748 42638 30880 42644
rect 30760 42622 30880 42638
rect 30760 42294 30788 42622
rect 31128 42566 31156 44814
rect 31208 44192 31260 44198
rect 31208 44134 31260 44140
rect 31220 43994 31248 44134
rect 31208 43988 31260 43994
rect 31208 43930 31260 43936
rect 31760 43172 31812 43178
rect 31760 43114 31812 43120
rect 31772 42770 31800 43114
rect 31760 42764 31812 42770
rect 31760 42706 31812 42712
rect 31116 42560 31168 42566
rect 31116 42502 31168 42508
rect 31760 42560 31812 42566
rect 31760 42502 31812 42508
rect 31024 42356 31076 42362
rect 31024 42298 31076 42304
rect 30748 42288 30800 42294
rect 30748 42230 30800 42236
rect 30656 41540 30708 41546
rect 30656 41482 30708 41488
rect 30668 41274 30696 41482
rect 30656 41268 30708 41274
rect 30656 41210 30708 41216
rect 30472 40044 30524 40050
rect 30472 39986 30524 39992
rect 30484 39642 30512 39986
rect 30564 39840 30616 39846
rect 30564 39782 30616 39788
rect 30472 39636 30524 39642
rect 30472 39578 30524 39584
rect 30576 39506 30604 39782
rect 30564 39500 30616 39506
rect 30564 39442 30616 39448
rect 30392 37726 30512 37754
rect 30380 37664 30432 37670
rect 30380 37606 30432 37612
rect 30392 37126 30420 37606
rect 30380 37120 30432 37126
rect 30380 37062 30432 37068
rect 30012 36916 30064 36922
rect 30012 36858 30064 36864
rect 30196 36916 30248 36922
rect 30196 36858 30248 36864
rect 29828 36848 29880 36854
rect 29828 36790 29880 36796
rect 30196 36780 30248 36786
rect 30196 36722 30248 36728
rect 30208 36666 30236 36722
rect 29932 36638 30236 36666
rect 29932 36582 29960 36638
rect 30484 36582 30512 37726
rect 29920 36576 29972 36582
rect 29920 36518 29972 36524
rect 30472 36576 30524 36582
rect 30472 36518 30524 36524
rect 29920 36168 29972 36174
rect 29920 36110 29972 36116
rect 29932 35290 29960 36110
rect 30012 35488 30064 35494
rect 30012 35430 30064 35436
rect 29920 35284 29972 35290
rect 29920 35226 29972 35232
rect 30024 35018 30052 35430
rect 30484 35222 30512 36518
rect 30760 35698 30788 42230
rect 31036 41750 31064 42298
rect 31128 42226 31156 42502
rect 31772 42294 31800 42502
rect 31760 42288 31812 42294
rect 31760 42230 31812 42236
rect 31116 42220 31168 42226
rect 31116 42162 31168 42168
rect 31024 41744 31076 41750
rect 31024 41686 31076 41692
rect 31300 41472 31352 41478
rect 31300 41414 31352 41420
rect 31956 41414 31984 63174
rect 32956 62824 33008 62830
rect 32956 62766 33008 62772
rect 33140 62824 33192 62830
rect 33140 62766 33192 62772
rect 32496 62756 32548 62762
rect 32496 62698 32548 62704
rect 32404 61192 32456 61198
rect 32404 61134 32456 61140
rect 32416 60110 32444 61134
rect 32404 60104 32456 60110
rect 32404 60046 32456 60052
rect 32220 60036 32272 60042
rect 32220 59978 32272 59984
rect 32232 59770 32260 59978
rect 32220 59764 32272 59770
rect 32220 59706 32272 59712
rect 32128 57860 32180 57866
rect 32128 57802 32180 57808
rect 32140 57526 32168 57802
rect 32128 57520 32180 57526
rect 32128 57462 32180 57468
rect 32312 56160 32364 56166
rect 32312 56102 32364 56108
rect 32324 55758 32352 56102
rect 32312 55752 32364 55758
rect 32312 55694 32364 55700
rect 32508 55282 32536 62698
rect 32968 61402 32996 62766
rect 33152 62490 33180 62766
rect 33140 62484 33192 62490
rect 33140 62426 33192 62432
rect 33428 61742 33456 63854
rect 34716 63578 34744 63922
rect 35348 63776 35400 63782
rect 35348 63718 35400 63724
rect 34934 63676 35242 63696
rect 34934 63674 34940 63676
rect 34996 63674 35020 63676
rect 35076 63674 35100 63676
rect 35156 63674 35180 63676
rect 35236 63674 35242 63676
rect 34996 63622 34998 63674
rect 35178 63622 35180 63674
rect 34934 63620 34940 63622
rect 34996 63620 35020 63622
rect 35076 63620 35100 63622
rect 35156 63620 35180 63622
rect 35236 63620 35242 63622
rect 34934 63600 35242 63620
rect 34704 63572 34756 63578
rect 34704 63514 34756 63520
rect 35360 63442 35388 63718
rect 35808 63572 35860 63578
rect 35808 63514 35860 63520
rect 36084 63572 36136 63578
rect 36084 63514 36136 63520
rect 35348 63436 35400 63442
rect 35348 63378 35400 63384
rect 35360 62966 35388 63378
rect 35716 63368 35768 63374
rect 35716 63310 35768 63316
rect 35348 62960 35400 62966
rect 35348 62902 35400 62908
rect 35440 62960 35492 62966
rect 35440 62902 35492 62908
rect 35452 62812 35480 62902
rect 35360 62784 35480 62812
rect 34934 62588 35242 62608
rect 34934 62586 34940 62588
rect 34996 62586 35020 62588
rect 35076 62586 35100 62588
rect 35156 62586 35180 62588
rect 35236 62586 35242 62588
rect 34996 62534 34998 62586
rect 35178 62534 35180 62586
rect 34934 62532 34940 62534
rect 34996 62532 35020 62534
rect 35076 62532 35100 62534
rect 35156 62532 35180 62534
rect 35236 62532 35242 62534
rect 34934 62512 35242 62532
rect 35360 62286 35388 62784
rect 35728 62762 35756 63310
rect 35716 62756 35768 62762
rect 35716 62698 35768 62704
rect 35440 62688 35492 62694
rect 35440 62630 35492 62636
rect 35452 62354 35480 62630
rect 35440 62348 35492 62354
rect 35440 62290 35492 62296
rect 34704 62280 34756 62286
rect 34704 62222 34756 62228
rect 35348 62280 35400 62286
rect 35348 62222 35400 62228
rect 33692 62144 33744 62150
rect 33692 62086 33744 62092
rect 33416 61736 33468 61742
rect 33416 61678 33468 61684
rect 33428 61402 33456 61678
rect 32956 61396 33008 61402
rect 32956 61338 33008 61344
rect 33416 61396 33468 61402
rect 33416 61338 33468 61344
rect 33704 60722 33732 62086
rect 34716 61606 34744 62222
rect 34796 61804 34848 61810
rect 34796 61746 34848 61752
rect 34704 61600 34756 61606
rect 34704 61542 34756 61548
rect 34716 61198 34744 61542
rect 34808 61334 34836 61746
rect 34934 61500 35242 61520
rect 34934 61498 34940 61500
rect 34996 61498 35020 61500
rect 35076 61498 35100 61500
rect 35156 61498 35180 61500
rect 35236 61498 35242 61500
rect 34996 61446 34998 61498
rect 35178 61446 35180 61498
rect 34934 61444 34940 61446
rect 34996 61444 35020 61446
rect 35076 61444 35100 61446
rect 35156 61444 35180 61446
rect 35236 61444 35242 61446
rect 34934 61424 35242 61444
rect 34796 61328 34848 61334
rect 34796 61270 34848 61276
rect 35360 61198 35388 62222
rect 35532 62144 35584 62150
rect 35532 62086 35584 62092
rect 34704 61192 34756 61198
rect 34704 61134 34756 61140
rect 35072 61192 35124 61198
rect 35072 61134 35124 61140
rect 35348 61192 35400 61198
rect 35348 61134 35400 61140
rect 33692 60716 33744 60722
rect 33692 60658 33744 60664
rect 33048 60036 33100 60042
rect 33048 59978 33100 59984
rect 32680 59628 32732 59634
rect 32680 59570 32732 59576
rect 32864 59628 32916 59634
rect 32864 59570 32916 59576
rect 32692 59226 32720 59570
rect 32680 59220 32732 59226
rect 32680 59162 32732 59168
rect 32588 58336 32640 58342
rect 32588 58278 32640 58284
rect 32600 57458 32628 58278
rect 32876 57458 32904 59570
rect 33060 57934 33088 59978
rect 33704 58546 33732 60658
rect 35084 60586 35112 61134
rect 35544 61130 35572 62086
rect 35820 61742 35848 63514
rect 36096 63238 36124 63514
rect 36084 63232 36136 63238
rect 36084 63174 36136 63180
rect 36280 62830 36308 65010
rect 36372 64598 36400 65010
rect 36544 65000 36596 65006
rect 36544 64942 36596 64948
rect 36360 64592 36412 64598
rect 36360 64534 36412 64540
rect 36556 64394 36584 64942
rect 36728 64592 36780 64598
rect 36728 64534 36780 64540
rect 36636 64456 36688 64462
rect 36636 64398 36688 64404
rect 36544 64388 36596 64394
rect 36544 64330 36596 64336
rect 36452 63436 36504 63442
rect 36452 63378 36504 63384
rect 36464 62898 36492 63378
rect 36360 62892 36412 62898
rect 36360 62834 36412 62840
rect 36452 62892 36504 62898
rect 36452 62834 36504 62840
rect 36084 62824 36136 62830
rect 36268 62824 36320 62830
rect 36136 62772 36216 62778
rect 36084 62766 36216 62772
rect 36268 62766 36320 62772
rect 36096 62750 36216 62766
rect 36188 62694 36216 62750
rect 35992 62688 36044 62694
rect 35992 62630 36044 62636
rect 36176 62688 36228 62694
rect 36176 62630 36228 62636
rect 36004 62422 36032 62630
rect 35992 62416 36044 62422
rect 35992 62358 36044 62364
rect 35808 61736 35860 61742
rect 35808 61678 35860 61684
rect 36084 61736 36136 61742
rect 36084 61678 36136 61684
rect 35992 61668 36044 61674
rect 35992 61610 36044 61616
rect 36004 61198 36032 61610
rect 36096 61334 36124 61678
rect 36084 61328 36136 61334
rect 36084 61270 36136 61276
rect 35992 61192 36044 61198
rect 35992 61134 36044 61140
rect 35532 61124 35584 61130
rect 35532 61066 35584 61072
rect 36004 60654 36032 61134
rect 36096 60722 36124 61270
rect 36372 61198 36400 62834
rect 36464 61810 36492 62834
rect 36556 62336 36584 64330
rect 36648 63578 36676 64398
rect 36740 64122 36768 64534
rect 36728 64116 36780 64122
rect 36728 64058 36780 64064
rect 36820 63980 36872 63986
rect 36820 63922 36872 63928
rect 36636 63572 36688 63578
rect 36636 63514 36688 63520
rect 36832 63374 36860 63922
rect 36820 63368 36872 63374
rect 36820 63310 36872 63316
rect 36636 63300 36688 63306
rect 36636 63242 36688 63248
rect 36648 62762 36676 63242
rect 36636 62756 36688 62762
rect 36636 62698 36688 62704
rect 36636 62348 36688 62354
rect 36556 62308 36636 62336
rect 36636 62290 36688 62296
rect 36648 62218 36676 62290
rect 36636 62212 36688 62218
rect 36636 62154 36688 62160
rect 36452 61804 36504 61810
rect 36452 61746 36504 61752
rect 36176 61192 36228 61198
rect 36176 61134 36228 61140
rect 36360 61192 36412 61198
rect 36360 61134 36412 61140
rect 36084 60716 36136 60722
rect 36084 60658 36136 60664
rect 35992 60648 36044 60654
rect 35992 60590 36044 60596
rect 35072 60580 35124 60586
rect 35072 60522 35124 60528
rect 33968 60512 34020 60518
rect 33968 60454 34020 60460
rect 33784 59968 33836 59974
rect 33784 59910 33836 59916
rect 33796 59634 33824 59910
rect 33980 59702 34008 60454
rect 34934 60412 35242 60432
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60336 35242 60356
rect 35348 59968 35400 59974
rect 35348 59910 35400 59916
rect 33968 59696 34020 59702
rect 33968 59638 34020 59644
rect 33784 59628 33836 59634
rect 33784 59570 33836 59576
rect 34934 59324 35242 59344
rect 34934 59322 34940 59324
rect 34996 59322 35020 59324
rect 35076 59322 35100 59324
rect 35156 59322 35180 59324
rect 35236 59322 35242 59324
rect 34996 59270 34998 59322
rect 35178 59270 35180 59322
rect 34934 59268 34940 59270
rect 34996 59268 35020 59270
rect 35076 59268 35100 59270
rect 35156 59268 35180 59270
rect 35236 59268 35242 59270
rect 34934 59248 35242 59268
rect 35360 58954 35388 59910
rect 36004 59566 36032 60590
rect 35992 59560 36044 59566
rect 35992 59502 36044 59508
rect 35348 58948 35400 58954
rect 35348 58890 35400 58896
rect 35348 58608 35400 58614
rect 35348 58550 35400 58556
rect 33692 58540 33744 58546
rect 33692 58482 33744 58488
rect 33876 58336 33928 58342
rect 33876 58278 33928 58284
rect 33048 57928 33100 57934
rect 33048 57870 33100 57876
rect 33060 57594 33088 57870
rect 33692 57792 33744 57798
rect 33692 57734 33744 57740
rect 33048 57588 33100 57594
rect 33048 57530 33100 57536
rect 32588 57452 32640 57458
rect 32588 57394 32640 57400
rect 32864 57452 32916 57458
rect 32864 57394 32916 57400
rect 33060 56302 33088 57530
rect 33704 57458 33732 57734
rect 33888 57526 33916 58278
rect 34934 58236 35242 58256
rect 34934 58234 34940 58236
rect 34996 58234 35020 58236
rect 35076 58234 35100 58236
rect 35156 58234 35180 58236
rect 35236 58234 35242 58236
rect 34996 58182 34998 58234
rect 35178 58182 35180 58234
rect 34934 58180 34940 58182
rect 34996 58180 35020 58182
rect 35076 58180 35100 58182
rect 35156 58180 35180 58182
rect 35236 58180 35242 58182
rect 34934 58160 35242 58180
rect 33968 57860 34020 57866
rect 33968 57802 34020 57808
rect 33876 57520 33928 57526
rect 33876 57462 33928 57468
rect 33692 57452 33744 57458
rect 33692 57394 33744 57400
rect 33980 57050 34008 57802
rect 34520 57384 34572 57390
rect 34520 57326 34572 57332
rect 34152 57248 34204 57254
rect 34152 57190 34204 57196
rect 33968 57044 34020 57050
rect 33968 56986 34020 56992
rect 34164 56846 34192 57190
rect 34152 56840 34204 56846
rect 34152 56782 34204 56788
rect 33324 56704 33376 56710
rect 33324 56646 33376 56652
rect 33336 56438 33364 56646
rect 33324 56432 33376 56438
rect 33324 56374 33376 56380
rect 33048 56296 33100 56302
rect 33048 56238 33100 56244
rect 32680 55684 32732 55690
rect 32680 55626 32732 55632
rect 32692 55418 32720 55626
rect 32680 55412 32732 55418
rect 32680 55354 32732 55360
rect 33060 55282 33088 56238
rect 34152 55684 34204 55690
rect 34152 55626 34204 55632
rect 32220 55276 32272 55282
rect 32220 55218 32272 55224
rect 32496 55276 32548 55282
rect 32496 55218 32548 55224
rect 33048 55276 33100 55282
rect 33048 55218 33100 55224
rect 32128 52352 32180 52358
rect 32128 52294 32180 52300
rect 32140 52086 32168 52294
rect 32128 52080 32180 52086
rect 32128 52022 32180 52028
rect 32036 51400 32088 51406
rect 32036 51342 32088 51348
rect 32048 49842 32076 51342
rect 32140 51338 32168 52022
rect 32128 51332 32180 51338
rect 32128 51274 32180 51280
rect 32036 49836 32088 49842
rect 32036 49778 32088 49784
rect 32036 46912 32088 46918
rect 32036 46854 32088 46860
rect 32048 46034 32076 46854
rect 32036 46028 32088 46034
rect 32036 45970 32088 45976
rect 32128 44192 32180 44198
rect 32128 44134 32180 44140
rect 32140 43790 32168 44134
rect 32128 43784 32180 43790
rect 32128 43726 32180 43732
rect 32128 42356 32180 42362
rect 32128 42298 32180 42304
rect 32140 42022 32168 42298
rect 32128 42016 32180 42022
rect 32128 41958 32180 41964
rect 31312 41070 31340 41414
rect 31956 41386 32076 41414
rect 31300 41064 31352 41070
rect 31300 41006 31352 41012
rect 31392 39840 31444 39846
rect 31392 39782 31444 39788
rect 31404 39438 31432 39782
rect 31024 39432 31076 39438
rect 31024 39374 31076 39380
rect 31392 39432 31444 39438
rect 31392 39374 31444 39380
rect 31036 39098 31064 39374
rect 31024 39092 31076 39098
rect 31024 39034 31076 39040
rect 30840 38956 30892 38962
rect 30840 38898 30892 38904
rect 30852 38350 30880 38898
rect 30840 38344 30892 38350
rect 30840 38286 30892 38292
rect 30852 36242 30880 38286
rect 31392 36712 31444 36718
rect 31392 36654 31444 36660
rect 30840 36236 30892 36242
rect 30840 36178 30892 36184
rect 30748 35692 30800 35698
rect 30748 35634 30800 35640
rect 30472 35216 30524 35222
rect 30472 35158 30524 35164
rect 30852 35086 30880 36178
rect 31300 36100 31352 36106
rect 31300 36042 31352 36048
rect 31312 35290 31340 36042
rect 31404 35698 31432 36654
rect 31392 35692 31444 35698
rect 31392 35634 31444 35640
rect 31300 35284 31352 35290
rect 31300 35226 31352 35232
rect 30840 35080 30892 35086
rect 30840 35022 30892 35028
rect 30012 35012 30064 35018
rect 30012 34954 30064 34960
rect 29736 34944 29788 34950
rect 29736 34886 29788 34892
rect 30196 34944 30248 34950
rect 30196 34886 30248 34892
rect 28816 34672 28868 34678
rect 28816 34614 28868 34620
rect 28828 32842 28856 34614
rect 28908 33992 28960 33998
rect 28908 33934 28960 33940
rect 29644 33992 29696 33998
rect 29644 33934 29696 33940
rect 28920 33454 28948 33934
rect 28908 33448 28960 33454
rect 28908 33390 28960 33396
rect 29656 32910 29684 33934
rect 29644 32904 29696 32910
rect 29644 32846 29696 32852
rect 28816 32836 28868 32842
rect 28816 32778 28868 32784
rect 29552 32768 29604 32774
rect 29552 32710 29604 32716
rect 29564 32502 29592 32710
rect 29644 32564 29696 32570
rect 29644 32506 29696 32512
rect 29552 32496 29604 32502
rect 29552 32438 29604 32444
rect 28724 32360 28776 32366
rect 28724 32302 28776 32308
rect 28736 32026 28764 32302
rect 28724 32020 28776 32026
rect 28724 31962 28776 31968
rect 29092 32020 29144 32026
rect 29092 31962 29144 31968
rect 28908 31884 28960 31890
rect 28908 31826 28960 31832
rect 28816 28960 28868 28966
rect 28816 28902 28868 28908
rect 28828 28150 28856 28902
rect 28816 28144 28868 28150
rect 28816 28086 28868 28092
rect 28828 27538 28856 28086
rect 28920 28014 28948 31826
rect 29000 29504 29052 29510
rect 29000 29446 29052 29452
rect 29012 29306 29040 29446
rect 29000 29300 29052 29306
rect 29000 29242 29052 29248
rect 29104 28762 29132 31962
rect 29656 31754 29684 32506
rect 29748 31890 29776 34886
rect 30208 34610 30236 34886
rect 30196 34604 30248 34610
rect 30196 34546 30248 34552
rect 30852 34202 30880 35022
rect 30472 34196 30524 34202
rect 30472 34138 30524 34144
rect 30840 34196 30892 34202
rect 30840 34138 30892 34144
rect 30104 33652 30156 33658
rect 30104 33594 30156 33600
rect 29828 33312 29880 33318
rect 29828 33254 29880 33260
rect 29736 31884 29788 31890
rect 29736 31826 29788 31832
rect 29644 31748 29696 31754
rect 29644 31690 29696 31696
rect 29736 31748 29788 31754
rect 29736 31690 29788 31696
rect 29644 30592 29696 30598
rect 29644 30534 29696 30540
rect 29656 30258 29684 30534
rect 29644 30252 29696 30258
rect 29644 30194 29696 30200
rect 29644 29640 29696 29646
rect 29644 29582 29696 29588
rect 29656 29306 29684 29582
rect 29644 29300 29696 29306
rect 29644 29242 29696 29248
rect 29644 29164 29696 29170
rect 29644 29106 29696 29112
rect 29092 28756 29144 28762
rect 29092 28698 29144 28704
rect 28908 28008 28960 28014
rect 28908 27950 28960 27956
rect 29104 27946 29132 28698
rect 29656 28558 29684 29106
rect 29644 28552 29696 28558
rect 29644 28494 29696 28500
rect 29748 28150 29776 31690
rect 29840 30122 29868 33254
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 29932 32026 29960 32846
rect 30116 32570 30144 33594
rect 30484 33522 30512 34138
rect 31404 33998 31432 35634
rect 31484 35488 31536 35494
rect 31484 35430 31536 35436
rect 31496 35086 31524 35430
rect 31576 35284 31628 35290
rect 31576 35226 31628 35232
rect 31484 35080 31536 35086
rect 31484 35022 31536 35028
rect 31588 34746 31616 35226
rect 31576 34740 31628 34746
rect 31576 34682 31628 34688
rect 31588 34066 31616 34682
rect 31576 34060 31628 34066
rect 31576 34002 31628 34008
rect 31392 33992 31444 33998
rect 31392 33934 31444 33940
rect 30472 33516 30524 33522
rect 30472 33458 30524 33464
rect 30564 33312 30616 33318
rect 30564 33254 30616 33260
rect 30104 32564 30156 32570
rect 30104 32506 30156 32512
rect 29920 32020 29972 32026
rect 29920 31962 29972 31968
rect 30576 31890 30604 33254
rect 31404 33130 31432 33934
rect 31312 33102 31432 33130
rect 30840 32768 30892 32774
rect 30840 32710 30892 32716
rect 30564 31884 30616 31890
rect 30564 31826 30616 31832
rect 30852 31822 30880 32710
rect 31312 32434 31340 33102
rect 31392 32904 31444 32910
rect 31392 32846 31444 32852
rect 31404 32570 31432 32846
rect 31392 32564 31444 32570
rect 31392 32506 31444 32512
rect 31300 32428 31352 32434
rect 31300 32370 31352 32376
rect 31852 32428 31904 32434
rect 31852 32370 31904 32376
rect 30840 31816 30892 31822
rect 30840 31758 30892 31764
rect 31392 31136 31444 31142
rect 31392 31078 31444 31084
rect 30472 30932 30524 30938
rect 30472 30874 30524 30880
rect 29828 30116 29880 30122
rect 29828 30058 29880 30064
rect 29840 29646 29868 30058
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29840 29102 29868 29582
rect 30288 29572 30340 29578
rect 30288 29514 30340 29520
rect 30300 29306 30328 29514
rect 30288 29300 30340 29306
rect 30288 29242 30340 29248
rect 29828 29096 29880 29102
rect 29828 29038 29880 29044
rect 30196 28416 30248 28422
rect 30196 28358 30248 28364
rect 29736 28144 29788 28150
rect 29736 28086 29788 28092
rect 30208 28082 30236 28358
rect 30196 28076 30248 28082
rect 30196 28018 30248 28024
rect 29092 27940 29144 27946
rect 29092 27882 29144 27888
rect 29184 27872 29236 27878
rect 29184 27814 29236 27820
rect 28816 27532 28868 27538
rect 28816 27474 28868 27480
rect 29196 27470 29224 27814
rect 30012 27532 30064 27538
rect 30012 27474 30064 27480
rect 29184 27464 29236 27470
rect 29184 27406 29236 27412
rect 28724 27328 28776 27334
rect 28724 27270 28776 27276
rect 28908 27328 28960 27334
rect 28908 27270 28960 27276
rect 29736 27328 29788 27334
rect 29736 27270 29788 27276
rect 28736 27130 28764 27270
rect 28724 27124 28776 27130
rect 28724 27066 28776 27072
rect 28920 26994 28948 27270
rect 29748 27062 29776 27270
rect 30024 27130 30052 27474
rect 30484 27470 30512 30874
rect 31404 30734 31432 31078
rect 31116 30728 31168 30734
rect 31116 30670 31168 30676
rect 31392 30728 31444 30734
rect 31392 30670 31444 30676
rect 31128 30394 31156 30670
rect 31760 30660 31812 30666
rect 31760 30602 31812 30608
rect 31116 30388 31168 30394
rect 31116 30330 31168 30336
rect 31772 30258 31800 30602
rect 31760 30252 31812 30258
rect 31760 30194 31812 30200
rect 31864 29646 31892 32370
rect 31944 32360 31996 32366
rect 31944 32302 31996 32308
rect 31956 31958 31984 32302
rect 31944 31952 31996 31958
rect 31944 31894 31996 31900
rect 31852 29640 31904 29646
rect 31852 29582 31904 29588
rect 31760 28620 31812 28626
rect 31760 28562 31812 28568
rect 31392 28416 31444 28422
rect 31392 28358 31444 28364
rect 31668 28416 31720 28422
rect 31668 28358 31720 28364
rect 31208 28076 31260 28082
rect 31208 28018 31260 28024
rect 31220 27674 31248 28018
rect 31208 27668 31260 27674
rect 31208 27610 31260 27616
rect 31404 27470 31432 28358
rect 31680 28218 31708 28358
rect 31668 28212 31720 28218
rect 31668 28154 31720 28160
rect 31772 27946 31800 28562
rect 31864 28558 31892 29582
rect 31944 29504 31996 29510
rect 31944 29446 31996 29452
rect 31956 29170 31984 29446
rect 31944 29164 31996 29170
rect 31944 29106 31996 29112
rect 31852 28552 31904 28558
rect 31852 28494 31904 28500
rect 31760 27940 31812 27946
rect 31760 27882 31812 27888
rect 30472 27464 30524 27470
rect 30472 27406 30524 27412
rect 31392 27464 31444 27470
rect 31392 27406 31444 27412
rect 30656 27328 30708 27334
rect 30656 27270 30708 27276
rect 30012 27124 30064 27130
rect 30012 27066 30064 27072
rect 29736 27056 29788 27062
rect 29736 26998 29788 27004
rect 30668 26994 30696 27270
rect 28908 26988 28960 26994
rect 28908 26930 28960 26936
rect 30656 26988 30708 26994
rect 30656 26930 30708 26936
rect 26436 26206 26648 26234
rect 28644 26206 28764 26234
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 25412 2576 25464 2582
rect 25412 2518 25464 2524
rect 25964 2576 26016 2582
rect 25964 2518 26016 2524
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 26620 2038 26648 26206
rect 28736 18358 28764 26206
rect 30668 25974 30696 26930
rect 31116 26376 31168 26382
rect 31116 26318 31168 26324
rect 31128 26042 31156 26318
rect 31116 26036 31168 26042
rect 31116 25978 31168 25984
rect 30656 25968 30708 25974
rect 30656 25910 30708 25916
rect 31392 25968 31444 25974
rect 31392 25910 31444 25916
rect 31404 24818 31432 25910
rect 31392 24812 31444 24818
rect 31392 24754 31444 24760
rect 32048 22094 32076 41386
rect 32128 38276 32180 38282
rect 32128 38218 32180 38224
rect 32140 38010 32168 38218
rect 32232 38214 32260 55218
rect 33324 54800 33376 54806
rect 33324 54742 33376 54748
rect 32404 54596 32456 54602
rect 32404 54538 32456 54544
rect 32416 53582 32444 54538
rect 33140 54324 33192 54330
rect 33140 54266 33192 54272
rect 32864 54188 32916 54194
rect 32864 54130 32916 54136
rect 32772 53984 32824 53990
rect 32772 53926 32824 53932
rect 32404 53576 32456 53582
rect 32404 53518 32456 53524
rect 32496 53100 32548 53106
rect 32496 53042 32548 53048
rect 32508 51882 32536 53042
rect 32784 53038 32812 53926
rect 32876 53786 32904 54130
rect 32864 53780 32916 53786
rect 32864 53722 32916 53728
rect 33152 53582 33180 54266
rect 33336 53582 33364 54742
rect 33140 53576 33192 53582
rect 33140 53518 33192 53524
rect 33324 53576 33376 53582
rect 33324 53518 33376 53524
rect 33416 53100 33468 53106
rect 33416 53042 33468 53048
rect 32772 53032 32824 53038
rect 32772 52974 32824 52980
rect 32680 52964 32732 52970
rect 32680 52906 32732 52912
rect 32496 51876 32548 51882
rect 32496 51818 32548 51824
rect 32496 50516 32548 50522
rect 32496 50458 32548 50464
rect 32508 48074 32536 50458
rect 32588 50312 32640 50318
rect 32588 50254 32640 50260
rect 32600 49978 32628 50254
rect 32588 49972 32640 49978
rect 32588 49914 32640 49920
rect 32600 49230 32628 49914
rect 32588 49224 32640 49230
rect 32588 49166 32640 49172
rect 32692 49162 32720 52906
rect 32784 51406 32812 52974
rect 33428 52698 33456 53042
rect 33416 52692 33468 52698
rect 33416 52634 33468 52640
rect 34164 52426 34192 55626
rect 34428 53508 34480 53514
rect 34428 53450 34480 53456
rect 34152 52420 34204 52426
rect 34152 52362 34204 52368
rect 34440 51474 34468 53450
rect 34428 51468 34480 51474
rect 34428 51410 34480 51416
rect 32772 51400 32824 51406
rect 32772 51342 32824 51348
rect 34152 51264 34204 51270
rect 34152 51206 34204 51212
rect 34164 50930 34192 51206
rect 34440 51074 34468 51410
rect 34348 51046 34468 51074
rect 34152 50924 34204 50930
rect 34152 50866 34204 50872
rect 34244 50788 34296 50794
rect 34244 50730 34296 50736
rect 33324 50176 33376 50182
rect 33324 50118 33376 50124
rect 32680 49156 32732 49162
rect 32680 49098 32732 49104
rect 33048 49156 33100 49162
rect 33048 49098 33100 49104
rect 32680 48272 32732 48278
rect 32680 48214 32732 48220
rect 32864 48272 32916 48278
rect 32956 48272 33008 48278
rect 32864 48214 32916 48220
rect 32954 48240 32956 48249
rect 33008 48240 33010 48249
rect 32692 48142 32720 48214
rect 32680 48136 32732 48142
rect 32680 48078 32732 48084
rect 32496 48068 32548 48074
rect 32496 48010 32548 48016
rect 32876 47666 32904 48214
rect 32954 48175 33010 48184
rect 32956 48000 33008 48006
rect 32956 47942 33008 47948
rect 32864 47660 32916 47666
rect 32864 47602 32916 47608
rect 32968 47258 32996 47942
rect 32956 47252 33008 47258
rect 32956 47194 33008 47200
rect 32496 47048 32548 47054
rect 32496 46990 32548 46996
rect 32508 46510 32536 46990
rect 32968 46714 32996 47194
rect 32956 46708 33008 46714
rect 32956 46650 33008 46656
rect 32496 46504 32548 46510
rect 32496 46446 32548 46452
rect 32772 46504 32824 46510
rect 32772 46446 32824 46452
rect 32864 46504 32916 46510
rect 32864 46446 32916 46452
rect 32508 44878 32536 46446
rect 32680 45824 32732 45830
rect 32680 45766 32732 45772
rect 32692 45558 32720 45766
rect 32680 45552 32732 45558
rect 32680 45494 32732 45500
rect 32496 44872 32548 44878
rect 32496 44814 32548 44820
rect 32496 42628 32548 42634
rect 32496 42570 32548 42576
rect 32508 42022 32536 42570
rect 32496 42016 32548 42022
rect 32496 41958 32548 41964
rect 32508 41138 32536 41958
rect 32692 41138 32720 45494
rect 32784 45098 32812 46446
rect 32876 45286 32904 46446
rect 32864 45280 32916 45286
rect 32864 45222 32916 45228
rect 32784 45070 32904 45098
rect 32772 43784 32824 43790
rect 32772 43726 32824 43732
rect 32784 43450 32812 43726
rect 32772 43444 32824 43450
rect 32772 43386 32824 43392
rect 32772 42832 32824 42838
rect 32772 42774 32824 42780
rect 32784 42702 32812 42774
rect 32772 42696 32824 42702
rect 32772 42638 32824 42644
rect 32772 42220 32824 42226
rect 32772 42162 32824 42168
rect 32784 41614 32812 42162
rect 32772 41608 32824 41614
rect 32772 41550 32824 41556
rect 32772 41472 32824 41478
rect 32772 41414 32824 41420
rect 32876 41414 32904 45070
rect 32956 43104 33008 43110
rect 32956 43046 33008 43052
rect 32968 42226 32996 43046
rect 32956 42220 33008 42226
rect 32956 42162 33008 42168
rect 32496 41132 32548 41138
rect 32496 41074 32548 41080
rect 32680 41132 32732 41138
rect 32680 41074 32732 41080
rect 32312 40044 32364 40050
rect 32312 39986 32364 39992
rect 32324 38962 32352 39986
rect 32680 39976 32732 39982
rect 32680 39918 32732 39924
rect 32692 39642 32720 39918
rect 32680 39636 32732 39642
rect 32680 39578 32732 39584
rect 32312 38956 32364 38962
rect 32312 38898 32364 38904
rect 32312 38752 32364 38758
rect 32312 38694 32364 38700
rect 32220 38208 32272 38214
rect 32220 38150 32272 38156
rect 32128 38004 32180 38010
rect 32128 37946 32180 37952
rect 32324 37874 32352 38694
rect 32312 37868 32364 37874
rect 32312 37810 32364 37816
rect 32680 37868 32732 37874
rect 32680 37810 32732 37816
rect 32692 36854 32720 37810
rect 32784 37262 32812 41414
rect 32876 41386 32996 41414
rect 32864 38752 32916 38758
rect 32864 38694 32916 38700
rect 32876 38554 32904 38694
rect 32864 38548 32916 38554
rect 32864 38490 32916 38496
rect 32772 37256 32824 37262
rect 32772 37198 32824 37204
rect 32680 36848 32732 36854
rect 32680 36790 32732 36796
rect 32968 36802 32996 41386
rect 33060 40526 33088 49098
rect 33140 48136 33192 48142
rect 33140 48078 33192 48084
rect 33152 47666 33180 48078
rect 33232 48068 33284 48074
rect 33232 48010 33284 48016
rect 33244 47977 33272 48010
rect 33230 47968 33286 47977
rect 33230 47903 33286 47912
rect 33140 47660 33192 47666
rect 33140 47602 33192 47608
rect 33048 40520 33100 40526
rect 33048 40462 33100 40468
rect 33232 40044 33284 40050
rect 33232 39986 33284 39992
rect 33244 39914 33272 39986
rect 33232 39908 33284 39914
rect 33232 39850 33284 39856
rect 33336 37874 33364 50118
rect 34256 49842 34284 50730
rect 34244 49836 34296 49842
rect 34244 49778 34296 49784
rect 33508 49632 33560 49638
rect 33508 49574 33560 49580
rect 33416 49156 33468 49162
rect 33416 49098 33468 49104
rect 33428 48550 33456 49098
rect 33520 49094 33548 49574
rect 33508 49088 33560 49094
rect 33508 49030 33560 49036
rect 33416 48544 33468 48550
rect 33416 48486 33468 48492
rect 33428 46578 33456 48486
rect 33520 46986 33548 49030
rect 33966 48240 34022 48249
rect 33692 48204 33744 48210
rect 33966 48175 33968 48184
rect 33692 48146 33744 48152
rect 34020 48175 34022 48184
rect 33968 48146 34020 48152
rect 33704 47598 33732 48146
rect 33876 48068 33928 48074
rect 33876 48010 33928 48016
rect 33888 47977 33916 48010
rect 33874 47968 33930 47977
rect 33874 47903 33930 47912
rect 33782 47832 33838 47841
rect 33782 47767 33784 47776
rect 33836 47767 33838 47776
rect 33968 47796 34020 47802
rect 33784 47738 33836 47744
rect 33968 47738 34020 47744
rect 33784 47660 33836 47666
rect 33784 47602 33836 47608
rect 33692 47592 33744 47598
rect 33692 47534 33744 47540
rect 33600 47456 33652 47462
rect 33600 47398 33652 47404
rect 33612 47122 33640 47398
rect 33600 47116 33652 47122
rect 33600 47058 33652 47064
rect 33508 46980 33560 46986
rect 33508 46922 33560 46928
rect 33416 46572 33468 46578
rect 33416 46514 33468 46520
rect 33520 46170 33548 46922
rect 33508 46164 33560 46170
rect 33508 46106 33560 46112
rect 33612 43738 33640 47058
rect 33796 46986 33824 47602
rect 33980 47258 34008 47738
rect 34348 47598 34376 51046
rect 34428 50856 34480 50862
rect 34428 50798 34480 50804
rect 34440 50250 34468 50798
rect 34428 50244 34480 50250
rect 34428 50186 34480 50192
rect 34440 48142 34468 50186
rect 34428 48136 34480 48142
rect 34428 48078 34480 48084
rect 34336 47592 34388 47598
rect 34336 47534 34388 47540
rect 33968 47252 34020 47258
rect 33968 47194 34020 47200
rect 34348 47122 34376 47534
rect 34336 47116 34388 47122
rect 34336 47058 34388 47064
rect 33784 46980 33836 46986
rect 33784 46922 33836 46928
rect 33796 46442 33824 46922
rect 33784 46436 33836 46442
rect 33784 46378 33836 46384
rect 34060 45960 34112 45966
rect 34060 45902 34112 45908
rect 34072 45354 34100 45902
rect 34532 45778 34560 57326
rect 34934 57148 35242 57168
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57072 35242 57092
rect 35360 56982 35388 58550
rect 36084 57792 36136 57798
rect 36084 57734 36136 57740
rect 36096 57458 36124 57734
rect 36084 57452 36136 57458
rect 36084 57394 36136 57400
rect 35900 57316 35952 57322
rect 35900 57258 35952 57264
rect 34796 56976 34848 56982
rect 34796 56918 34848 56924
rect 35348 56976 35400 56982
rect 35348 56918 35400 56924
rect 34612 56228 34664 56234
rect 34612 56170 34664 56176
rect 34624 55894 34652 56170
rect 34612 55888 34664 55894
rect 34612 55830 34664 55836
rect 34808 55826 34836 56918
rect 35072 56772 35124 56778
rect 35072 56714 35124 56720
rect 35348 56772 35400 56778
rect 35348 56714 35400 56720
rect 35084 56506 35112 56714
rect 35072 56500 35124 56506
rect 35072 56442 35124 56448
rect 34934 56060 35242 56080
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55984 35242 56004
rect 34796 55820 34848 55826
rect 34796 55762 34848 55768
rect 34612 55616 34664 55622
rect 34612 55558 34664 55564
rect 34624 49337 34652 55558
rect 34704 55276 34756 55282
rect 34704 55218 34756 55224
rect 34716 54874 34744 55218
rect 34934 54972 35242 54992
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54896 35242 54916
rect 34704 54868 34756 54874
rect 34704 54810 34756 54816
rect 34934 53884 35242 53904
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53808 35242 53828
rect 35256 53576 35308 53582
rect 35256 53518 35308 53524
rect 35268 53242 35296 53518
rect 34796 53236 34848 53242
rect 34796 53178 34848 53184
rect 35256 53236 35308 53242
rect 35256 53178 35308 53184
rect 34808 52086 34836 53178
rect 34934 52796 35242 52816
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52720 35242 52740
rect 34796 52080 34848 52086
rect 34796 52022 34848 52028
rect 34934 51708 35242 51728
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51632 35242 51652
rect 34888 51536 34940 51542
rect 34888 51478 34940 51484
rect 34900 51406 34928 51478
rect 34704 51400 34756 51406
rect 34704 51342 34756 51348
rect 34888 51400 34940 51406
rect 34888 51342 34940 51348
rect 34716 50998 34744 51342
rect 34704 50992 34756 50998
rect 34704 50934 34756 50940
rect 34934 50620 35242 50640
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50544 35242 50564
rect 34796 49632 34848 49638
rect 34796 49574 34848 49580
rect 34610 49328 34666 49337
rect 34610 49263 34666 49272
rect 34704 49224 34756 49230
rect 34704 49166 34756 49172
rect 34612 49156 34664 49162
rect 34612 49098 34664 49104
rect 34624 48890 34652 49098
rect 34612 48884 34664 48890
rect 34612 48826 34664 48832
rect 34716 48686 34744 49166
rect 34808 48754 34836 49574
rect 34934 49532 35242 49552
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49456 35242 49476
rect 34886 49328 34942 49337
rect 34886 49263 34942 49272
rect 34796 48748 34848 48754
rect 34796 48690 34848 48696
rect 34704 48680 34756 48686
rect 34900 48634 34928 49263
rect 34704 48622 34756 48628
rect 34716 47734 34744 48622
rect 34808 48606 34928 48634
rect 34704 47728 34756 47734
rect 34704 47670 34756 47676
rect 34612 47456 34664 47462
rect 34612 47398 34664 47404
rect 34624 45898 34652 47398
rect 34612 45892 34664 45898
rect 34612 45834 34664 45840
rect 34532 45750 34652 45778
rect 34520 45552 34572 45558
rect 34520 45494 34572 45500
rect 34428 45416 34480 45422
rect 34428 45358 34480 45364
rect 34060 45348 34112 45354
rect 34060 45290 34112 45296
rect 34336 44736 34388 44742
rect 34336 44678 34388 44684
rect 34152 44396 34204 44402
rect 34152 44338 34204 44344
rect 33784 44192 33836 44198
rect 33784 44134 33836 44140
rect 33796 43790 33824 44134
rect 33784 43784 33836 43790
rect 33612 43710 33732 43738
rect 33784 43726 33836 43732
rect 33600 43648 33652 43654
rect 33600 43590 33652 43596
rect 33612 43382 33640 43590
rect 33600 43376 33652 43382
rect 33600 43318 33652 43324
rect 33416 42152 33468 42158
rect 33416 42094 33468 42100
rect 33428 38962 33456 42094
rect 33508 41064 33560 41070
rect 33508 41006 33560 41012
rect 33520 40458 33548 41006
rect 33508 40452 33560 40458
rect 33508 40394 33560 40400
rect 33612 39914 33640 43318
rect 33704 41414 33732 43710
rect 34164 43450 34192 44338
rect 34152 43444 34204 43450
rect 34152 43386 34204 43392
rect 33968 43376 34020 43382
rect 33968 43318 34020 43324
rect 33876 43308 33928 43314
rect 33876 43250 33928 43256
rect 33784 42628 33836 42634
rect 33784 42570 33836 42576
rect 33796 42158 33824 42570
rect 33888 42208 33916 43250
rect 33980 42566 34008 43318
rect 34152 42696 34204 42702
rect 34152 42638 34204 42644
rect 33968 42560 34020 42566
rect 33968 42502 34020 42508
rect 34164 42362 34192 42638
rect 34152 42356 34204 42362
rect 34152 42298 34204 42304
rect 33968 42220 34020 42226
rect 33888 42180 33968 42208
rect 33968 42162 34020 42168
rect 33784 42152 33836 42158
rect 33784 42094 33836 42100
rect 33980 41614 34008 42162
rect 33968 41608 34020 41614
rect 33968 41550 34020 41556
rect 34348 41414 34376 44678
rect 34440 43994 34468 45358
rect 34532 44418 34560 45494
rect 34624 44538 34652 45750
rect 34716 45558 34744 47670
rect 34808 47462 34836 48606
rect 34934 48444 35242 48464
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48368 35242 48388
rect 34796 47456 34848 47462
rect 34796 47398 34848 47404
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 34796 47184 34848 47190
rect 34796 47126 34848 47132
rect 34808 45966 34836 47126
rect 35360 46510 35388 56714
rect 35912 56166 35940 57258
rect 35992 56296 36044 56302
rect 35992 56238 36044 56244
rect 35808 56160 35860 56166
rect 35808 56102 35860 56108
rect 35900 56160 35952 56166
rect 35900 56102 35952 56108
rect 35820 55842 35848 56102
rect 35820 55814 35940 55842
rect 35912 55690 35940 55814
rect 35900 55684 35952 55690
rect 35900 55626 35952 55632
rect 35532 55276 35584 55282
rect 35532 55218 35584 55224
rect 35440 55072 35492 55078
rect 35440 55014 35492 55020
rect 35452 54670 35480 55014
rect 35440 54664 35492 54670
rect 35440 54606 35492 54612
rect 35440 53644 35492 53650
rect 35440 53586 35492 53592
rect 35452 52426 35480 53586
rect 35544 53174 35572 55218
rect 36004 55146 36032 56238
rect 36096 55826 36124 57394
rect 36188 57322 36216 61134
rect 36372 60858 36400 61134
rect 36544 61056 36596 61062
rect 36544 60998 36596 61004
rect 36360 60852 36412 60858
rect 36360 60794 36412 60800
rect 36556 60722 36584 60998
rect 36544 60716 36596 60722
rect 36544 60658 36596 60664
rect 36544 60104 36596 60110
rect 36544 60046 36596 60052
rect 36556 59770 36584 60046
rect 36544 59764 36596 59770
rect 36544 59706 36596 59712
rect 36268 59560 36320 59566
rect 36268 59502 36320 59508
rect 36280 59226 36308 59502
rect 36648 59498 36676 62154
rect 36360 59492 36412 59498
rect 36360 59434 36412 59440
rect 36636 59492 36688 59498
rect 36636 59434 36688 59440
rect 36268 59220 36320 59226
rect 36268 59162 36320 59168
rect 36268 57928 36320 57934
rect 36268 57870 36320 57876
rect 36280 57594 36308 57870
rect 36268 57588 36320 57594
rect 36268 57530 36320 57536
rect 36176 57316 36228 57322
rect 36176 57258 36228 57264
rect 36280 56914 36308 57530
rect 36268 56908 36320 56914
rect 36268 56850 36320 56856
rect 36176 56364 36228 56370
rect 36176 56306 36228 56312
rect 36084 55820 36136 55826
rect 36084 55762 36136 55768
rect 36096 55282 36124 55762
rect 36084 55276 36136 55282
rect 36084 55218 36136 55224
rect 35992 55140 36044 55146
rect 35992 55082 36044 55088
rect 35808 55072 35860 55078
rect 35808 55014 35860 55020
rect 35716 54868 35768 54874
rect 35716 54810 35768 54816
rect 35728 54754 35756 54810
rect 35636 54726 35756 54754
rect 35636 53582 35664 54726
rect 35716 54664 35768 54670
rect 35716 54606 35768 54612
rect 35624 53576 35676 53582
rect 35624 53518 35676 53524
rect 35728 53514 35756 54606
rect 35716 53508 35768 53514
rect 35716 53450 35768 53456
rect 35532 53168 35584 53174
rect 35532 53110 35584 53116
rect 35728 53106 35756 53450
rect 35716 53100 35768 53106
rect 35636 53060 35716 53088
rect 35532 52964 35584 52970
rect 35532 52906 35584 52912
rect 35544 52630 35572 52906
rect 35532 52624 35584 52630
rect 35532 52566 35584 52572
rect 35440 52420 35492 52426
rect 35440 52362 35492 52368
rect 35544 51882 35572 52566
rect 35532 51876 35584 51882
rect 35532 51818 35584 51824
rect 35636 51814 35664 53060
rect 35716 53042 35768 53048
rect 35716 52896 35768 52902
rect 35716 52838 35768 52844
rect 35624 51808 35676 51814
rect 35624 51750 35676 51756
rect 35624 51400 35676 51406
rect 35624 51342 35676 51348
rect 35532 51264 35584 51270
rect 35532 51206 35584 51212
rect 35544 51074 35572 51206
rect 35452 51046 35572 51074
rect 35452 50998 35480 51046
rect 35440 50992 35492 50998
rect 35440 50934 35492 50940
rect 35452 49842 35480 50934
rect 35636 50708 35664 51342
rect 35728 51270 35756 52838
rect 35820 51406 35848 55014
rect 35992 53576 36044 53582
rect 35992 53518 36044 53524
rect 35900 53440 35952 53446
rect 35900 53382 35952 53388
rect 35912 53242 35940 53382
rect 35900 53236 35952 53242
rect 35900 53178 35952 53184
rect 36004 52086 36032 53518
rect 36084 53032 36136 53038
rect 36084 52974 36136 52980
rect 35992 52080 36044 52086
rect 35992 52022 36044 52028
rect 36004 51542 36032 52022
rect 35992 51536 36044 51542
rect 35992 51478 36044 51484
rect 35808 51400 35860 51406
rect 35808 51342 35860 51348
rect 35716 51264 35768 51270
rect 35716 51206 35768 51212
rect 35820 50998 35848 51342
rect 36096 51338 36124 52974
rect 36084 51332 36136 51338
rect 36084 51274 36136 51280
rect 35808 50992 35860 50998
rect 35808 50934 35860 50940
rect 35716 50720 35768 50726
rect 35544 50680 35716 50708
rect 35544 49842 35572 50680
rect 35716 50662 35768 50668
rect 35716 50176 35768 50182
rect 35716 50118 35768 50124
rect 35440 49836 35492 49842
rect 35440 49778 35492 49784
rect 35532 49836 35584 49842
rect 35532 49778 35584 49784
rect 35452 49434 35480 49778
rect 35440 49428 35492 49434
rect 35440 49370 35492 49376
rect 35544 49314 35572 49778
rect 35452 49286 35572 49314
rect 35452 47802 35480 49286
rect 35624 48136 35676 48142
rect 35624 48078 35676 48084
rect 35440 47796 35492 47802
rect 35440 47738 35492 47744
rect 35532 47728 35584 47734
rect 35532 47670 35584 47676
rect 35440 47456 35492 47462
rect 35440 47398 35492 47404
rect 35452 47122 35480 47398
rect 35440 47116 35492 47122
rect 35440 47058 35492 47064
rect 35544 46986 35572 47670
rect 35636 47666 35664 48078
rect 35624 47660 35676 47666
rect 35624 47602 35676 47608
rect 35624 47524 35676 47530
rect 35624 47466 35676 47472
rect 35532 46980 35584 46986
rect 35532 46922 35584 46928
rect 35348 46504 35400 46510
rect 35348 46446 35400 46452
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 35544 45966 35572 46922
rect 35636 46714 35664 47466
rect 35624 46708 35676 46714
rect 35624 46650 35676 46656
rect 34796 45960 34848 45966
rect 34796 45902 34848 45908
rect 35532 45960 35584 45966
rect 35532 45902 35584 45908
rect 34704 45552 34756 45558
rect 34704 45494 34756 45500
rect 34716 44946 34744 45494
rect 34808 45422 34836 45902
rect 35624 45824 35676 45830
rect 35624 45766 35676 45772
rect 35636 45490 35664 45766
rect 35624 45484 35676 45490
rect 35624 45426 35676 45432
rect 34796 45416 34848 45422
rect 34796 45358 34848 45364
rect 35728 45354 35756 50118
rect 35820 49842 35848 50934
rect 36084 50312 36136 50318
rect 36084 50254 36136 50260
rect 36096 49910 36124 50254
rect 36084 49904 36136 49910
rect 36084 49846 36136 49852
rect 35808 49836 35860 49842
rect 35808 49778 35860 49784
rect 36188 48142 36216 56306
rect 36268 55752 36320 55758
rect 36268 55694 36320 55700
rect 36280 55350 36308 55694
rect 36268 55344 36320 55350
rect 36268 55286 36320 55292
rect 36268 55140 36320 55146
rect 36268 55082 36320 55088
rect 36176 48136 36228 48142
rect 36176 48078 36228 48084
rect 35990 47832 36046 47841
rect 35808 47796 35860 47802
rect 35990 47767 35992 47776
rect 35808 47738 35860 47744
rect 36044 47767 36046 47776
rect 35992 47738 36044 47744
rect 35820 47122 35848 47738
rect 35808 47116 35860 47122
rect 35808 47058 35860 47064
rect 35900 46572 35952 46578
rect 35900 46514 35952 46520
rect 35716 45348 35768 45354
rect 35716 45290 35768 45296
rect 35440 45280 35492 45286
rect 35440 45222 35492 45228
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34704 44940 34756 44946
rect 34704 44882 34756 44888
rect 34716 44538 34744 44882
rect 35452 44878 35480 45222
rect 35440 44872 35492 44878
rect 35440 44814 35492 44820
rect 34612 44532 34664 44538
rect 34612 44474 34664 44480
rect 34704 44532 34756 44538
rect 34704 44474 34756 44480
rect 34532 44390 34744 44418
rect 34520 44328 34572 44334
rect 34520 44270 34572 44276
rect 34612 44328 34664 44334
rect 34612 44270 34664 44276
rect 34428 43988 34480 43994
rect 34428 43930 34480 43936
rect 34440 43110 34468 43930
rect 34532 43858 34560 44270
rect 34520 43852 34572 43858
rect 34520 43794 34572 43800
rect 34532 43382 34560 43794
rect 34520 43376 34572 43382
rect 34520 43318 34572 43324
rect 34428 43104 34480 43110
rect 34428 43046 34480 43052
rect 34520 43104 34572 43110
rect 34520 43046 34572 43052
rect 34440 42906 34468 43046
rect 34428 42900 34480 42906
rect 34428 42842 34480 42848
rect 33704 41386 33824 41414
rect 34348 41386 34468 41414
rect 33600 39908 33652 39914
rect 33600 39850 33652 39856
rect 33600 39364 33652 39370
rect 33600 39306 33652 39312
rect 33416 38956 33468 38962
rect 33416 38898 33468 38904
rect 33612 38894 33640 39306
rect 33600 38888 33652 38894
rect 33600 38830 33652 38836
rect 33796 38282 33824 41386
rect 34440 41138 34468 41386
rect 34428 41132 34480 41138
rect 34428 41074 34480 41080
rect 34532 41070 34560 43046
rect 34520 41064 34572 41070
rect 34520 41006 34572 41012
rect 33876 40928 33928 40934
rect 33876 40870 33928 40876
rect 33888 39914 33916 40870
rect 34532 40730 34560 41006
rect 34520 40724 34572 40730
rect 34520 40666 34572 40672
rect 34244 39976 34296 39982
rect 34244 39918 34296 39924
rect 33876 39908 33928 39914
rect 33876 39850 33928 39856
rect 33888 38826 33916 39850
rect 34256 39642 34284 39918
rect 34244 39636 34296 39642
rect 34244 39578 34296 39584
rect 34428 38888 34480 38894
rect 34428 38830 34480 38836
rect 33876 38820 33928 38826
rect 33876 38762 33928 38768
rect 34060 38820 34112 38826
rect 34060 38762 34112 38768
rect 34072 38282 34100 38762
rect 34440 38758 34468 38830
rect 34428 38752 34480 38758
rect 34428 38694 34480 38700
rect 33784 38276 33836 38282
rect 33784 38218 33836 38224
rect 34060 38276 34112 38282
rect 34060 38218 34112 38224
rect 34520 38276 34572 38282
rect 34520 38218 34572 38224
rect 33324 37868 33376 37874
rect 33324 37810 33376 37816
rect 33232 37800 33284 37806
rect 33232 37742 33284 37748
rect 32968 36774 33088 36802
rect 32310 36680 32366 36689
rect 32310 36615 32366 36624
rect 32324 36378 32352 36615
rect 32312 36372 32364 36378
rect 32312 36314 32364 36320
rect 32324 35766 32352 36314
rect 32312 35760 32364 35766
rect 32312 35702 32364 35708
rect 32404 35692 32456 35698
rect 32404 35634 32456 35640
rect 32312 34604 32364 34610
rect 32312 34546 32364 34552
rect 32324 34202 32352 34546
rect 32312 34196 32364 34202
rect 32312 34138 32364 34144
rect 32416 33810 32444 35634
rect 32588 35488 32640 35494
rect 32588 35430 32640 35436
rect 32600 35154 32628 35430
rect 32588 35148 32640 35154
rect 32588 35090 32640 35096
rect 32324 33782 32444 33810
rect 32324 32434 32352 33782
rect 33060 33454 33088 36774
rect 33244 36378 33272 37742
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 33324 36780 33376 36786
rect 33324 36722 33376 36728
rect 33232 36372 33284 36378
rect 33232 36314 33284 36320
rect 33140 35488 33192 35494
rect 33140 35430 33192 35436
rect 33152 35086 33180 35430
rect 33140 35080 33192 35086
rect 33140 35022 33192 35028
rect 33244 34932 33272 36314
rect 33336 36038 33364 36722
rect 33520 36378 33548 37198
rect 33508 36372 33560 36378
rect 33508 36314 33560 36320
rect 33324 36032 33376 36038
rect 33324 35974 33376 35980
rect 33152 34904 33272 34932
rect 33152 34406 33180 34904
rect 33336 34762 33364 35974
rect 33416 35692 33468 35698
rect 33416 35634 33468 35640
rect 33244 34734 33364 34762
rect 33428 34746 33456 35634
rect 33416 34740 33468 34746
rect 33244 34678 33272 34734
rect 33416 34682 33468 34688
rect 33232 34672 33284 34678
rect 33232 34614 33284 34620
rect 33140 34400 33192 34406
rect 33140 34342 33192 34348
rect 33048 33448 33100 33454
rect 33048 33390 33100 33396
rect 33152 33318 33180 34342
rect 33244 33590 33272 34614
rect 33796 34134 33824 38218
rect 33876 37120 33928 37126
rect 33876 37062 33928 37068
rect 33888 36786 33916 37062
rect 33876 36780 33928 36786
rect 33876 36722 33928 36728
rect 33888 36106 33916 36722
rect 34532 36650 34560 38218
rect 34520 36644 34572 36650
rect 34520 36586 34572 36592
rect 33876 36100 33928 36106
rect 33876 36042 33928 36048
rect 34532 35222 34560 36586
rect 34520 35216 34572 35222
rect 34520 35158 34572 35164
rect 33968 35080 34020 35086
rect 33968 35022 34020 35028
rect 33980 34950 34008 35022
rect 33968 34944 34020 34950
rect 33968 34886 34020 34892
rect 33980 34610 34008 34886
rect 33968 34604 34020 34610
rect 33968 34546 34020 34552
rect 33784 34128 33836 34134
rect 33784 34070 33836 34076
rect 34060 33856 34112 33862
rect 34060 33798 34112 33804
rect 33232 33584 33284 33590
rect 33232 33526 33284 33532
rect 33140 33312 33192 33318
rect 33140 33254 33192 33260
rect 32404 32904 32456 32910
rect 32404 32846 32456 32852
rect 32416 32570 32444 32846
rect 32864 32836 32916 32842
rect 32864 32778 32916 32784
rect 32404 32564 32456 32570
rect 32404 32506 32456 32512
rect 32312 32428 32364 32434
rect 32312 32370 32364 32376
rect 32324 31346 32352 32370
rect 32876 32026 32904 32778
rect 32956 32292 33008 32298
rect 32956 32234 33008 32240
rect 32864 32020 32916 32026
rect 32864 31962 32916 31968
rect 32220 31340 32272 31346
rect 32220 31282 32272 31288
rect 32312 31340 32364 31346
rect 32312 31282 32364 31288
rect 32232 30394 32260 31282
rect 32324 30666 32352 31282
rect 32312 30660 32364 30666
rect 32312 30602 32364 30608
rect 32496 30592 32548 30598
rect 32496 30534 32548 30540
rect 32220 30388 32272 30394
rect 32220 30330 32272 30336
rect 32508 30326 32536 30534
rect 32128 30320 32180 30326
rect 32128 30262 32180 30268
rect 32496 30320 32548 30326
rect 32496 30262 32548 30268
rect 32140 29170 32168 30262
rect 32680 30116 32732 30122
rect 32680 30058 32732 30064
rect 32692 29782 32720 30058
rect 32680 29776 32732 29782
rect 32680 29718 32732 29724
rect 32128 29164 32180 29170
rect 32128 29106 32180 29112
rect 32496 29096 32548 29102
rect 32496 29038 32548 29044
rect 32128 26308 32180 26314
rect 32128 26250 32180 26256
rect 32140 26042 32168 26250
rect 32128 26036 32180 26042
rect 32128 25978 32180 25984
rect 32508 25362 32536 29038
rect 32680 27464 32732 27470
rect 32680 27406 32732 27412
rect 32692 27130 32720 27406
rect 32864 27328 32916 27334
rect 32864 27270 32916 27276
rect 32680 27124 32732 27130
rect 32680 27066 32732 27072
rect 32876 26382 32904 27270
rect 32968 26450 32996 32234
rect 33152 30938 33180 33254
rect 33140 30932 33192 30938
rect 33140 30874 33192 30880
rect 33244 30802 33272 33526
rect 33784 33516 33836 33522
rect 33784 33458 33836 33464
rect 33324 33312 33376 33318
rect 33324 33254 33376 33260
rect 33336 31822 33364 33254
rect 33796 33114 33824 33458
rect 33784 33108 33836 33114
rect 33784 33050 33836 33056
rect 33600 32836 33652 32842
rect 33600 32778 33652 32784
rect 33612 32366 33640 32778
rect 33796 32434 33824 33050
rect 33784 32428 33836 32434
rect 33784 32370 33836 32376
rect 33600 32360 33652 32366
rect 33600 32302 33652 32308
rect 34072 32298 34100 33798
rect 34428 32360 34480 32366
rect 34428 32302 34480 32308
rect 34060 32292 34112 32298
rect 34060 32234 34112 32240
rect 33968 31884 34020 31890
rect 33968 31826 34020 31832
rect 33324 31816 33376 31822
rect 33324 31758 33376 31764
rect 33324 31136 33376 31142
rect 33324 31078 33376 31084
rect 33232 30796 33284 30802
rect 33232 30738 33284 30744
rect 33244 30326 33272 30738
rect 33336 30666 33364 31078
rect 33416 30932 33468 30938
rect 33416 30874 33468 30880
rect 33324 30660 33376 30666
rect 33324 30602 33376 30608
rect 33232 30320 33284 30326
rect 33232 30262 33284 30268
rect 33336 30258 33364 30602
rect 33324 30252 33376 30258
rect 33324 30194 33376 30200
rect 33428 30122 33456 30874
rect 33416 30116 33468 30122
rect 33416 30058 33468 30064
rect 33980 29306 34008 31826
rect 34072 31754 34100 32234
rect 34440 31958 34468 32302
rect 34428 31952 34480 31958
rect 34428 31894 34480 31900
rect 34072 31726 34192 31754
rect 34060 30184 34112 30190
rect 34060 30126 34112 30132
rect 33968 29300 34020 29306
rect 33968 29242 34020 29248
rect 33140 29096 33192 29102
rect 33060 29044 33140 29050
rect 33060 29038 33192 29044
rect 33060 29022 33180 29038
rect 33060 28626 33088 29022
rect 33048 28620 33100 28626
rect 33048 28562 33100 28568
rect 33232 27872 33284 27878
rect 33232 27814 33284 27820
rect 33244 27470 33272 27814
rect 34072 27606 34100 30126
rect 34164 30122 34192 31726
rect 34520 31408 34572 31414
rect 34520 31350 34572 31356
rect 34532 30598 34560 31350
rect 34520 30592 34572 30598
rect 34520 30534 34572 30540
rect 34532 30394 34560 30534
rect 34520 30388 34572 30394
rect 34520 30330 34572 30336
rect 34520 30184 34572 30190
rect 34520 30126 34572 30132
rect 34152 30116 34204 30122
rect 34152 30058 34204 30064
rect 34164 29034 34192 30058
rect 34428 30048 34480 30054
rect 34428 29990 34480 29996
rect 34440 29850 34468 29990
rect 34428 29844 34480 29850
rect 34428 29786 34480 29792
rect 34532 29714 34560 30126
rect 34520 29708 34572 29714
rect 34520 29650 34572 29656
rect 34152 29028 34204 29034
rect 34152 28970 34204 28976
rect 34336 28008 34388 28014
rect 34336 27950 34388 27956
rect 34520 28008 34572 28014
rect 34520 27950 34572 27956
rect 34060 27600 34112 27606
rect 34060 27542 34112 27548
rect 34348 27470 34376 27950
rect 34532 27538 34560 27950
rect 34520 27532 34572 27538
rect 34520 27474 34572 27480
rect 33232 27464 33284 27470
rect 33232 27406 33284 27412
rect 33968 27464 34020 27470
rect 33968 27406 34020 27412
rect 34336 27464 34388 27470
rect 34336 27406 34388 27412
rect 33980 26994 34008 27406
rect 34244 27396 34296 27402
rect 34244 27338 34296 27344
rect 34256 27062 34284 27338
rect 34244 27056 34296 27062
rect 34244 26998 34296 27004
rect 33140 26988 33192 26994
rect 33140 26930 33192 26936
rect 33968 26988 34020 26994
rect 33968 26930 34020 26936
rect 32956 26444 33008 26450
rect 32956 26386 33008 26392
rect 33152 26382 33180 26930
rect 32864 26376 32916 26382
rect 32864 26318 32916 26324
rect 33140 26376 33192 26382
rect 33140 26318 33192 26324
rect 33784 26376 33836 26382
rect 33784 26318 33836 26324
rect 32496 25356 32548 25362
rect 32496 25298 32548 25304
rect 32404 25152 32456 25158
rect 32404 25094 32456 25100
rect 32220 24812 32272 24818
rect 32220 24754 32272 24760
rect 32232 24410 32260 24754
rect 32220 24404 32272 24410
rect 32220 24346 32272 24352
rect 32416 24206 32444 25094
rect 32508 24614 32536 25298
rect 33152 25294 33180 26318
rect 33324 26240 33376 26246
rect 33324 26182 33376 26188
rect 33336 25906 33364 26182
rect 33796 25974 33824 26318
rect 33784 25968 33836 25974
rect 33784 25910 33836 25916
rect 33324 25900 33376 25906
rect 33324 25842 33376 25848
rect 33692 25832 33744 25838
rect 33692 25774 33744 25780
rect 33704 25498 33732 25774
rect 33692 25492 33744 25498
rect 33692 25434 33744 25440
rect 33796 25294 33824 25910
rect 33968 25900 34020 25906
rect 33968 25842 34020 25848
rect 33140 25288 33192 25294
rect 33140 25230 33192 25236
rect 33784 25288 33836 25294
rect 33784 25230 33836 25236
rect 33980 24954 34008 25842
rect 33968 24948 34020 24954
rect 33968 24890 34020 24896
rect 32496 24608 32548 24614
rect 32496 24550 32548 24556
rect 32404 24200 32456 24206
rect 32404 24142 32456 24148
rect 31956 22066 32076 22094
rect 28724 18352 28776 18358
rect 28724 18294 28776 18300
rect 27436 18216 27488 18222
rect 27436 18158 27488 18164
rect 27448 2514 27476 18158
rect 31956 12782 31984 22066
rect 32128 12844 32180 12850
rect 32128 12786 32180 12792
rect 31944 12776 31996 12782
rect 31944 12718 31996 12724
rect 27436 2508 27488 2514
rect 27436 2450 27488 2456
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 26608 2032 26660 2038
rect 26608 1974 26660 1980
rect 27080 800 27108 2382
rect 28368 800 28396 2382
rect 32140 2310 32168 12786
rect 32404 12640 32456 12646
rect 32404 12582 32456 12588
rect 32416 6914 32444 12582
rect 32324 6886 32444 6914
rect 32324 2650 32352 6886
rect 34624 4146 34652 44270
rect 34716 40390 34744 44390
rect 34796 44396 34848 44402
rect 34796 44338 34848 44344
rect 34808 42022 34836 44338
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 35808 43920 35860 43926
rect 35808 43862 35860 43868
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 35440 42628 35492 42634
rect 35440 42570 35492 42576
rect 35452 42362 35480 42570
rect 35716 42560 35768 42566
rect 35716 42502 35768 42508
rect 35440 42356 35492 42362
rect 35440 42298 35492 42304
rect 35532 42356 35584 42362
rect 35532 42298 35584 42304
rect 35544 42226 35572 42298
rect 35728 42226 35756 42502
rect 35532 42220 35584 42226
rect 35532 42162 35584 42168
rect 35716 42220 35768 42226
rect 35716 42162 35768 42168
rect 34796 42016 34848 42022
rect 34796 41958 34848 41964
rect 34808 41546 34836 41958
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 35440 41608 35492 41614
rect 35440 41550 35492 41556
rect 35532 41608 35584 41614
rect 35532 41550 35584 41556
rect 34796 41540 34848 41546
rect 34796 41482 34848 41488
rect 35256 41472 35308 41478
rect 35256 41414 35308 41420
rect 35268 41206 35296 41414
rect 35256 41200 35308 41206
rect 35256 41142 35308 41148
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 35452 40730 35480 41550
rect 35544 40934 35572 41550
rect 35532 40928 35584 40934
rect 35532 40870 35584 40876
rect 35624 40928 35676 40934
rect 35624 40870 35676 40876
rect 34796 40724 34848 40730
rect 34796 40666 34848 40672
rect 35348 40724 35400 40730
rect 35348 40666 35400 40672
rect 35440 40724 35492 40730
rect 35440 40666 35492 40672
rect 34704 40384 34756 40390
rect 34704 40326 34756 40332
rect 34808 39982 34836 40666
rect 35360 40474 35388 40666
rect 35164 40452 35216 40458
rect 35360 40446 35480 40474
rect 35636 40458 35664 40870
rect 35164 40394 35216 40400
rect 35176 40186 35204 40394
rect 35348 40384 35400 40390
rect 35348 40326 35400 40332
rect 35164 40180 35216 40186
rect 35164 40122 35216 40128
rect 34796 39976 34848 39982
rect 34796 39918 34848 39924
rect 34808 38894 34836 39918
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 35256 39364 35308 39370
rect 35256 39306 35308 39312
rect 35268 39098 35296 39306
rect 35360 39302 35388 40326
rect 35452 39642 35480 40446
rect 35624 40452 35676 40458
rect 35624 40394 35676 40400
rect 35440 39636 35492 39642
rect 35440 39578 35492 39584
rect 35452 39522 35480 39578
rect 35452 39494 35572 39522
rect 35440 39432 35492 39438
rect 35440 39374 35492 39380
rect 35348 39296 35400 39302
rect 35348 39238 35400 39244
rect 35256 39092 35308 39098
rect 35256 39034 35308 39040
rect 34796 38888 34848 38894
rect 34796 38830 34848 38836
rect 35348 38888 35400 38894
rect 35348 38830 35400 38836
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34704 37800 34756 37806
rect 34704 37742 34756 37748
rect 34716 36174 34744 37742
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34796 36712 34848 36718
rect 34888 36712 34940 36718
rect 34796 36654 34848 36660
rect 34886 36680 34888 36689
rect 35360 36700 35388 38830
rect 35452 38554 35480 39374
rect 35440 38548 35492 38554
rect 35440 38490 35492 38496
rect 35440 37732 35492 37738
rect 35440 37674 35492 37680
rect 35452 37330 35480 37674
rect 35440 37324 35492 37330
rect 35440 37266 35492 37272
rect 35440 36712 35492 36718
rect 34940 36680 34942 36689
rect 35360 36672 35440 36700
rect 34704 36168 34756 36174
rect 34704 36110 34756 36116
rect 34716 31686 34744 36110
rect 34704 31680 34756 31686
rect 34704 31622 34756 31628
rect 34704 31340 34756 31346
rect 34704 31282 34756 31288
rect 34716 30938 34744 31282
rect 34704 30932 34756 30938
rect 34704 30874 34756 30880
rect 34704 30184 34756 30190
rect 34704 30126 34756 30132
rect 34716 29782 34744 30126
rect 34704 29776 34756 29782
rect 34704 29718 34756 29724
rect 34716 29102 34744 29718
rect 34704 29096 34756 29102
rect 34704 29038 34756 29044
rect 34704 28960 34756 28966
rect 34704 28902 34756 28908
rect 34716 28762 34744 28902
rect 34704 28756 34756 28762
rect 34704 28698 34756 28704
rect 34808 28200 34836 36654
rect 35440 36654 35492 36660
rect 34886 36615 34942 36624
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 35452 36394 35480 36654
rect 35544 36582 35572 39494
rect 35820 38962 35848 43862
rect 35912 43178 35940 46514
rect 36188 46170 36216 48078
rect 36280 46714 36308 55082
rect 36372 51406 36400 59434
rect 36544 57792 36596 57798
rect 36544 57734 36596 57740
rect 36556 56846 36584 57734
rect 36544 56840 36596 56846
rect 36544 56782 36596 56788
rect 36728 56432 36780 56438
rect 36728 56374 36780 56380
rect 36636 56228 36688 56234
rect 36636 56170 36688 56176
rect 36648 55826 36676 56170
rect 36636 55820 36688 55826
rect 36636 55762 36688 55768
rect 36636 55616 36688 55622
rect 36636 55558 36688 55564
rect 36648 55418 36676 55558
rect 36636 55412 36688 55418
rect 36636 55354 36688 55360
rect 36740 55350 36768 56374
rect 36820 55956 36872 55962
rect 36820 55898 36872 55904
rect 36832 55758 36860 55898
rect 36820 55752 36872 55758
rect 36820 55694 36872 55700
rect 36728 55344 36780 55350
rect 36728 55286 36780 55292
rect 36740 54754 36768 55286
rect 36648 54726 36768 54754
rect 36648 52698 36676 54726
rect 36728 54596 36780 54602
rect 36728 54538 36780 54544
rect 36636 52692 36688 52698
rect 36556 52652 36636 52680
rect 36452 51536 36504 51542
rect 36452 51478 36504 51484
rect 36360 51400 36412 51406
rect 36360 51342 36412 51348
rect 36464 49774 36492 51478
rect 36556 50930 36584 52652
rect 36636 52634 36688 52640
rect 36740 51406 36768 54538
rect 36728 51400 36780 51406
rect 36728 51342 36780 51348
rect 36820 51060 36872 51066
rect 36820 51002 36872 51008
rect 36544 50924 36596 50930
rect 36544 50866 36596 50872
rect 36556 50318 36584 50866
rect 36636 50788 36688 50794
rect 36636 50730 36688 50736
rect 36544 50312 36596 50318
rect 36544 50254 36596 50260
rect 36648 50250 36676 50730
rect 36832 50522 36860 51002
rect 36820 50516 36872 50522
rect 36820 50458 36872 50464
rect 36636 50244 36688 50250
rect 36636 50186 36688 50192
rect 36544 49836 36596 49842
rect 36544 49778 36596 49784
rect 36452 49768 36504 49774
rect 36452 49710 36504 49716
rect 36556 49162 36584 49778
rect 36648 49230 36676 50186
rect 36636 49224 36688 49230
rect 36636 49166 36688 49172
rect 36544 49156 36596 49162
rect 36544 49098 36596 49104
rect 36358 48104 36414 48113
rect 36358 48039 36414 48048
rect 36372 47734 36400 48039
rect 36360 47728 36412 47734
rect 36360 47670 36412 47676
rect 36452 47048 36504 47054
rect 36452 46990 36504 46996
rect 36728 47048 36780 47054
rect 36728 46990 36780 46996
rect 36360 46980 36412 46986
rect 36360 46922 36412 46928
rect 36268 46708 36320 46714
rect 36268 46650 36320 46656
rect 36176 46164 36228 46170
rect 36176 46106 36228 46112
rect 36268 45280 36320 45286
rect 36268 45222 36320 45228
rect 36176 44736 36228 44742
rect 36176 44678 36228 44684
rect 36188 43858 36216 44678
rect 36280 44470 36308 45222
rect 36268 44464 36320 44470
rect 36268 44406 36320 44412
rect 36268 44192 36320 44198
rect 36268 44134 36320 44140
rect 36176 43852 36228 43858
rect 36176 43794 36228 43800
rect 36280 43790 36308 44134
rect 36372 43994 36400 46922
rect 36464 45898 36492 46990
rect 36740 46578 36768 46990
rect 36728 46572 36780 46578
rect 36728 46514 36780 46520
rect 36452 45892 36504 45898
rect 36452 45834 36504 45840
rect 36360 43988 36412 43994
rect 36360 43930 36412 43936
rect 36268 43784 36320 43790
rect 36268 43726 36320 43732
rect 35992 43716 36044 43722
rect 35992 43658 36044 43664
rect 35900 43172 35952 43178
rect 35900 43114 35952 43120
rect 36004 42226 36032 43658
rect 36280 42770 36308 43726
rect 36268 42764 36320 42770
rect 36268 42706 36320 42712
rect 36084 42560 36136 42566
rect 36084 42502 36136 42508
rect 35992 42220 36044 42226
rect 35992 42162 36044 42168
rect 36096 42158 36124 42502
rect 36084 42152 36136 42158
rect 36084 42094 36136 42100
rect 36464 41414 36492 45834
rect 36544 42220 36596 42226
rect 36544 42162 36596 42168
rect 36556 41546 36584 42162
rect 36544 41540 36596 41546
rect 36544 41482 36596 41488
rect 36280 41386 36492 41414
rect 35808 38956 35860 38962
rect 35808 38898 35860 38904
rect 35820 37874 35848 38898
rect 35992 38752 36044 38758
rect 35992 38694 36044 38700
rect 36004 38282 36032 38694
rect 35992 38276 36044 38282
rect 35992 38218 36044 38224
rect 35808 37868 35860 37874
rect 35808 37810 35860 37816
rect 36004 37330 36032 38218
rect 35624 37324 35676 37330
rect 35624 37266 35676 37272
rect 35992 37324 36044 37330
rect 35992 37266 36044 37272
rect 35532 36576 35584 36582
rect 35532 36518 35584 36524
rect 35452 36366 35572 36394
rect 35348 35556 35400 35562
rect 35348 35498 35400 35504
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 35256 35148 35308 35154
rect 35256 35090 35308 35096
rect 35268 34746 35296 35090
rect 35256 34740 35308 34746
rect 35256 34682 35308 34688
rect 35268 34490 35296 34682
rect 35360 34610 35388 35498
rect 35544 35494 35572 36366
rect 35636 35698 35664 37266
rect 35808 37256 35860 37262
rect 35808 37198 35860 37204
rect 35820 36786 35848 37198
rect 35992 37120 36044 37126
rect 35992 37062 36044 37068
rect 35808 36780 35860 36786
rect 35808 36722 35860 36728
rect 35716 36576 35768 36582
rect 35716 36518 35768 36524
rect 35624 35692 35676 35698
rect 35624 35634 35676 35640
rect 35440 35488 35492 35494
rect 35440 35430 35492 35436
rect 35532 35488 35584 35494
rect 35532 35430 35584 35436
rect 35452 34610 35480 35430
rect 35636 35193 35664 35634
rect 35622 35184 35678 35193
rect 35622 35119 35678 35128
rect 35624 35080 35676 35086
rect 35624 35022 35676 35028
rect 35636 34898 35664 35022
rect 35544 34870 35664 34898
rect 35348 34604 35400 34610
rect 35348 34546 35400 34552
rect 35440 34604 35492 34610
rect 35440 34546 35492 34552
rect 35268 34462 35388 34490
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 35360 33930 35388 34462
rect 35348 33924 35400 33930
rect 35348 33866 35400 33872
rect 35440 33448 35492 33454
rect 35440 33390 35492 33396
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34888 32768 34940 32774
rect 34888 32710 34940 32716
rect 34900 32570 34928 32710
rect 34888 32564 34940 32570
rect 34888 32506 34940 32512
rect 35452 32434 35480 33390
rect 35440 32428 35492 32434
rect 35440 32370 35492 32376
rect 35348 32360 35400 32366
rect 35348 32302 35400 32308
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 35360 30818 35388 32302
rect 35440 31408 35492 31414
rect 35440 31350 35492 31356
rect 34900 30790 35388 30818
rect 34900 30190 34928 30790
rect 35348 30660 35400 30666
rect 35348 30602 35400 30608
rect 34888 30184 34940 30190
rect 34888 30126 34940 30132
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 35360 29850 35388 30602
rect 35348 29844 35400 29850
rect 35348 29786 35400 29792
rect 35452 29730 35480 31350
rect 35268 29702 35480 29730
rect 35268 29306 35296 29702
rect 35256 29300 35308 29306
rect 35256 29242 35308 29248
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 35164 28552 35216 28558
rect 35164 28494 35216 28500
rect 35176 28218 35204 28494
rect 34716 28172 34836 28200
rect 35164 28212 35216 28218
rect 34716 27146 34744 28172
rect 35164 28154 35216 28160
rect 34796 28076 34848 28082
rect 34796 28018 34848 28024
rect 34808 27606 34836 28018
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34796 27600 34848 27606
rect 34796 27542 34848 27548
rect 34716 27118 34836 27146
rect 35544 27130 35572 34870
rect 35622 34776 35678 34785
rect 35622 34711 35678 34720
rect 35636 32994 35664 34711
rect 35728 34202 35756 36518
rect 35716 34196 35768 34202
rect 35716 34138 35768 34144
rect 35728 33522 35756 34138
rect 35820 33862 35848 36722
rect 36004 36242 36032 37062
rect 36176 36848 36228 36854
rect 36176 36790 36228 36796
rect 36188 36378 36216 36790
rect 36176 36372 36228 36378
rect 36176 36314 36228 36320
rect 35992 36236 36044 36242
rect 35992 36178 36044 36184
rect 36280 35850 36308 41386
rect 36728 39296 36780 39302
rect 36728 39238 36780 39244
rect 36740 38962 36768 39238
rect 36728 38956 36780 38962
rect 36728 38898 36780 38904
rect 36544 38752 36596 38758
rect 36544 38694 36596 38700
rect 36556 38350 36584 38694
rect 36544 38344 36596 38350
rect 36544 38286 36596 38292
rect 36544 36576 36596 36582
rect 36544 36518 36596 36524
rect 36360 36100 36412 36106
rect 36360 36042 36412 36048
rect 36188 35834 36308 35850
rect 36372 35834 36400 36042
rect 36176 35828 36308 35834
rect 36228 35822 36308 35828
rect 36360 35828 36412 35834
rect 36176 35770 36228 35776
rect 36360 35770 36412 35776
rect 36556 35698 36584 36518
rect 36544 35692 36596 35698
rect 36544 35634 36596 35640
rect 35992 35624 36044 35630
rect 35992 35566 36044 35572
rect 35900 35488 35952 35494
rect 35900 35430 35952 35436
rect 35912 35154 35940 35430
rect 35900 35148 35952 35154
rect 35900 35090 35952 35096
rect 36004 34202 36032 35566
rect 35992 34196 36044 34202
rect 35992 34138 36044 34144
rect 35808 33856 35860 33862
rect 35808 33798 35860 33804
rect 35716 33516 35768 33522
rect 35716 33458 35768 33464
rect 35728 33114 35756 33458
rect 35716 33108 35768 33114
rect 35716 33050 35768 33056
rect 35636 32966 35756 32994
rect 35624 32904 35676 32910
rect 35624 32846 35676 32852
rect 35636 32026 35664 32846
rect 35624 32020 35676 32026
rect 35624 31962 35676 31968
rect 35728 31822 35756 32966
rect 35820 32570 35848 33798
rect 36452 32836 36504 32842
rect 36452 32778 36504 32784
rect 36464 32570 36492 32778
rect 36636 32768 36688 32774
rect 36636 32710 36688 32716
rect 35808 32564 35860 32570
rect 35808 32506 35860 32512
rect 36452 32564 36504 32570
rect 36452 32506 36504 32512
rect 35716 31816 35768 31822
rect 35716 31758 35768 31764
rect 35624 31680 35676 31686
rect 35624 31622 35676 31628
rect 35636 28082 35664 31622
rect 35728 31346 35756 31758
rect 35820 31414 35848 32506
rect 36648 32434 36676 32710
rect 36636 32428 36688 32434
rect 36636 32370 36688 32376
rect 35900 32224 35952 32230
rect 35900 32166 35952 32172
rect 35912 31754 35940 32166
rect 35912 31726 36032 31754
rect 35808 31408 35860 31414
rect 35808 31350 35860 31356
rect 35716 31340 35768 31346
rect 35716 31282 35768 31288
rect 36004 31210 36032 31726
rect 35992 31204 36044 31210
rect 35992 31146 36044 31152
rect 35716 31136 35768 31142
rect 35716 31078 35768 31084
rect 35728 29646 35756 31078
rect 35716 29640 35768 29646
rect 35716 29582 35768 29588
rect 36004 29034 36032 31146
rect 36176 31136 36228 31142
rect 36176 31078 36228 31084
rect 36188 30734 36216 31078
rect 36176 30728 36228 30734
rect 36176 30670 36228 30676
rect 36544 29096 36596 29102
rect 36544 29038 36596 29044
rect 35992 29028 36044 29034
rect 35992 28970 36044 28976
rect 35900 28960 35952 28966
rect 35900 28902 35952 28908
rect 35912 28558 35940 28902
rect 36556 28762 36584 29038
rect 36544 28756 36596 28762
rect 36544 28698 36596 28704
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 35624 28076 35676 28082
rect 35624 28018 35676 28024
rect 34704 26988 34756 26994
rect 34704 26930 34756 26936
rect 34716 26586 34744 26930
rect 34704 26580 34756 26586
rect 34704 26522 34756 26528
rect 34808 26042 34836 27118
rect 35532 27124 35584 27130
rect 35532 27066 35584 27072
rect 35440 26988 35492 26994
rect 35440 26930 35492 26936
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 35452 26586 35480 26930
rect 35624 26784 35676 26790
rect 35624 26726 35676 26732
rect 35440 26580 35492 26586
rect 35440 26522 35492 26528
rect 35636 26382 35664 26726
rect 35624 26376 35676 26382
rect 35624 26318 35676 26324
rect 34796 26036 34848 26042
rect 34796 25978 34848 25984
rect 34808 25294 34836 25978
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34796 25288 34848 25294
rect 34796 25230 34848 25236
rect 35072 25152 35124 25158
rect 35072 25094 35124 25100
rect 35084 24818 35112 25094
rect 35072 24812 35124 24818
rect 35072 24754 35124 24760
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 36924 18086 36952 69226
rect 37280 69216 37332 69222
rect 37280 69158 37332 69164
rect 37292 68338 37320 69158
rect 37280 68332 37332 68338
rect 37280 68274 37332 68280
rect 38028 68270 38056 71200
rect 39028 69216 39080 69222
rect 39028 69158 39080 69164
rect 38936 68808 38988 68814
rect 38936 68750 38988 68756
rect 37556 68264 37608 68270
rect 37556 68206 37608 68212
rect 38016 68264 38068 68270
rect 38016 68206 38068 68212
rect 37568 67930 37596 68206
rect 37556 67924 37608 67930
rect 37556 67866 37608 67872
rect 37464 67720 37516 67726
rect 37464 67662 37516 67668
rect 37004 67108 37056 67114
rect 37004 67050 37056 67056
rect 37016 33046 37044 67050
rect 37476 66502 37504 67662
rect 38568 67652 38620 67658
rect 38568 67594 38620 67600
rect 37464 66496 37516 66502
rect 37464 66438 37516 66444
rect 38292 65068 38344 65074
rect 38292 65010 38344 65016
rect 38200 64864 38252 64870
rect 38200 64806 38252 64812
rect 38212 64462 38240 64806
rect 38304 64666 38332 65010
rect 38292 64660 38344 64666
rect 38292 64602 38344 64608
rect 38200 64456 38252 64462
rect 38200 64398 38252 64404
rect 38108 64388 38160 64394
rect 38108 64330 38160 64336
rect 37280 64320 37332 64326
rect 37280 64262 37332 64268
rect 37740 64320 37792 64326
rect 37740 64262 37792 64268
rect 37292 64122 37320 64262
rect 37280 64116 37332 64122
rect 37280 64058 37332 64064
rect 37648 64048 37700 64054
rect 37648 63990 37700 63996
rect 37660 63918 37688 63990
rect 37752 63986 37780 64262
rect 38016 64116 38068 64122
rect 38016 64058 38068 64064
rect 37740 63980 37792 63986
rect 37740 63922 37792 63928
rect 37648 63912 37700 63918
rect 37648 63854 37700 63860
rect 37280 63776 37332 63782
rect 37280 63718 37332 63724
rect 37292 63442 37320 63718
rect 37280 63436 37332 63442
rect 37280 63378 37332 63384
rect 37660 62898 37688 63854
rect 38028 63442 38056 64058
rect 38016 63436 38068 63442
rect 38016 63378 38068 63384
rect 37740 63368 37792 63374
rect 37740 63310 37792 63316
rect 37648 62892 37700 62898
rect 37648 62834 37700 62840
rect 37660 62422 37688 62834
rect 37648 62416 37700 62422
rect 37648 62358 37700 62364
rect 37372 61192 37424 61198
rect 37372 61134 37424 61140
rect 37384 60734 37412 61134
rect 37292 60706 37412 60734
rect 37292 59566 37320 60706
rect 37372 59628 37424 59634
rect 37372 59570 37424 59576
rect 37280 59560 37332 59566
rect 37280 59502 37332 59508
rect 37292 59090 37320 59502
rect 37280 59084 37332 59090
rect 37280 59026 37332 59032
rect 37384 58682 37412 59570
rect 37464 58880 37516 58886
rect 37464 58822 37516 58828
rect 37372 58676 37424 58682
rect 37372 58618 37424 58624
rect 37476 58546 37504 58822
rect 37464 58540 37516 58546
rect 37464 58482 37516 58488
rect 37648 57928 37700 57934
rect 37648 57870 37700 57876
rect 37556 57588 37608 57594
rect 37556 57530 37608 57536
rect 37372 57452 37424 57458
rect 37372 57394 37424 57400
rect 37384 56506 37412 57394
rect 37372 56500 37424 56506
rect 37372 56442 37424 56448
rect 37384 56370 37412 56442
rect 37372 56364 37424 56370
rect 37372 56306 37424 56312
rect 37188 56296 37240 56302
rect 37188 56238 37240 56244
rect 37096 56160 37148 56166
rect 37096 56102 37148 56108
rect 37108 53242 37136 56102
rect 37200 55758 37228 56238
rect 37188 55752 37240 55758
rect 37188 55694 37240 55700
rect 37188 55616 37240 55622
rect 37188 55558 37240 55564
rect 37200 55282 37228 55558
rect 37188 55276 37240 55282
rect 37188 55218 37240 55224
rect 37096 53236 37148 53242
rect 37096 53178 37148 53184
rect 37108 51338 37136 53178
rect 37096 51332 37148 51338
rect 37096 51274 37148 51280
rect 37096 50516 37148 50522
rect 37096 50458 37148 50464
rect 37108 50182 37136 50458
rect 37096 50176 37148 50182
rect 37096 50118 37148 50124
rect 37108 49774 37136 50118
rect 37096 49768 37148 49774
rect 37096 49710 37148 49716
rect 37200 34474 37228 55218
rect 37280 53508 37332 53514
rect 37280 53450 37332 53456
rect 37292 53242 37320 53450
rect 37280 53236 37332 53242
rect 37280 53178 37332 53184
rect 37280 52624 37332 52630
rect 37280 52566 37332 52572
rect 37292 49638 37320 52566
rect 37384 49978 37412 56306
rect 37568 54194 37596 57530
rect 37660 57526 37688 57870
rect 37648 57520 37700 57526
rect 37648 57462 37700 57468
rect 37648 57384 37700 57390
rect 37648 57326 37700 57332
rect 37660 57050 37688 57326
rect 37648 57044 37700 57050
rect 37648 56986 37700 56992
rect 37556 54188 37608 54194
rect 37556 54130 37608 54136
rect 37464 53780 37516 53786
rect 37464 53722 37516 53728
rect 37476 53106 37504 53722
rect 37568 53582 37596 54130
rect 37556 53576 37608 53582
rect 37556 53518 37608 53524
rect 37464 53100 37516 53106
rect 37464 53042 37516 53048
rect 37476 52630 37504 53042
rect 37464 52624 37516 52630
rect 37464 52566 37516 52572
rect 37568 52018 37596 53518
rect 37556 52012 37608 52018
rect 37556 51954 37608 51960
rect 37648 51808 37700 51814
rect 37648 51750 37700 51756
rect 37660 51406 37688 51750
rect 37648 51400 37700 51406
rect 37648 51342 37700 51348
rect 37648 50448 37700 50454
rect 37648 50390 37700 50396
rect 37556 50244 37608 50250
rect 37556 50186 37608 50192
rect 37464 50176 37516 50182
rect 37464 50118 37516 50124
rect 37372 49972 37424 49978
rect 37372 49914 37424 49920
rect 37280 49632 37332 49638
rect 37280 49574 37332 49580
rect 37292 49094 37320 49574
rect 37280 49088 37332 49094
rect 37280 49030 37332 49036
rect 37384 48906 37412 49914
rect 37476 49756 37504 50118
rect 37568 49910 37596 50186
rect 37660 49978 37688 50390
rect 37752 50182 37780 63310
rect 37924 62892 37976 62898
rect 37924 62834 37976 62840
rect 37936 62490 37964 62834
rect 38028 62762 38056 63378
rect 38120 62830 38148 64330
rect 38108 62824 38160 62830
rect 38108 62766 38160 62772
rect 38016 62756 38068 62762
rect 38016 62698 38068 62704
rect 37924 62484 37976 62490
rect 37924 62426 37976 62432
rect 38028 62286 38056 62698
rect 38016 62280 38068 62286
rect 38016 62222 38068 62228
rect 38120 61198 38148 62766
rect 38200 62688 38252 62694
rect 38200 62630 38252 62636
rect 38212 62286 38240 62630
rect 38200 62280 38252 62286
rect 38200 62222 38252 62228
rect 38108 61192 38160 61198
rect 38108 61134 38160 61140
rect 38120 60722 38148 61134
rect 38108 60716 38160 60722
rect 38108 60658 38160 60664
rect 38016 58948 38068 58954
rect 38016 58890 38068 58896
rect 38028 58138 38056 58890
rect 38016 58132 38068 58138
rect 38016 58074 38068 58080
rect 37832 55072 37884 55078
rect 37832 55014 37884 55020
rect 37844 53990 37872 55014
rect 37832 53984 37884 53990
rect 37832 53926 37884 53932
rect 37844 53038 37872 53926
rect 37924 53440 37976 53446
rect 37924 53382 37976 53388
rect 37936 53174 37964 53382
rect 37924 53168 37976 53174
rect 37924 53110 37976 53116
rect 37832 53032 37884 53038
rect 37832 52974 37884 52980
rect 37924 52012 37976 52018
rect 37924 51954 37976 51960
rect 37936 51610 37964 51954
rect 37924 51604 37976 51610
rect 37924 51546 37976 51552
rect 38028 50794 38056 58074
rect 38200 56772 38252 56778
rect 38200 56714 38252 56720
rect 38212 56234 38240 56714
rect 38200 56228 38252 56234
rect 38200 56170 38252 56176
rect 38212 55758 38240 56170
rect 38200 55752 38252 55758
rect 38200 55694 38252 55700
rect 38108 54528 38160 54534
rect 38108 54470 38160 54476
rect 38292 54528 38344 54534
rect 38292 54470 38344 54476
rect 38016 50788 38068 50794
rect 38016 50730 38068 50736
rect 38028 50182 38056 50730
rect 37740 50176 37792 50182
rect 37740 50118 37792 50124
rect 38016 50176 38068 50182
rect 38016 50118 38068 50124
rect 37648 49972 37700 49978
rect 37648 49914 37700 49920
rect 37556 49904 37608 49910
rect 37556 49846 37608 49852
rect 37476 49728 37596 49756
rect 37464 49088 37516 49094
rect 37464 49030 37516 49036
rect 37292 48878 37412 48906
rect 37292 48142 37320 48878
rect 37372 48748 37424 48754
rect 37372 48690 37424 48696
rect 37384 48278 37412 48690
rect 37372 48272 37424 48278
rect 37372 48214 37424 48220
rect 37280 48136 37332 48142
rect 37280 48078 37332 48084
rect 37280 46980 37332 46986
rect 37280 46922 37332 46928
rect 37292 46578 37320 46922
rect 37280 46572 37332 46578
rect 37280 46514 37332 46520
rect 37476 45558 37504 49030
rect 37568 48550 37596 49728
rect 37648 49156 37700 49162
rect 37648 49098 37700 49104
rect 37556 48544 37608 48550
rect 37556 48486 37608 48492
rect 37464 45552 37516 45558
rect 37464 45494 37516 45500
rect 37556 45484 37608 45490
rect 37556 45426 37608 45432
rect 37464 45280 37516 45286
rect 37464 45222 37516 45228
rect 37372 42696 37424 42702
rect 37372 42638 37424 42644
rect 37384 42226 37412 42638
rect 37372 42220 37424 42226
rect 37372 42162 37424 42168
rect 37280 41744 37332 41750
rect 37278 41712 37280 41721
rect 37332 41712 37334 41721
rect 37278 41647 37334 41656
rect 37384 41562 37412 42162
rect 37292 41546 37412 41562
rect 37280 41540 37412 41546
rect 37332 41534 37412 41540
rect 37280 41482 37332 41488
rect 37280 41132 37332 41138
rect 37280 41074 37332 41080
rect 37292 40594 37320 41074
rect 37280 40588 37332 40594
rect 37280 40530 37332 40536
rect 37384 40526 37412 41534
rect 37476 41478 37504 45222
rect 37568 45082 37596 45426
rect 37556 45076 37608 45082
rect 37556 45018 37608 45024
rect 37660 42634 37688 49098
rect 37924 48544 37976 48550
rect 37924 48486 37976 48492
rect 37936 48074 37964 48486
rect 38120 48314 38148 54470
rect 38304 54262 38332 54470
rect 38292 54256 38344 54262
rect 38292 54198 38344 54204
rect 38476 50924 38528 50930
rect 38476 50866 38528 50872
rect 38488 50522 38516 50866
rect 38476 50516 38528 50522
rect 38476 50458 38528 50464
rect 38580 50318 38608 67594
rect 38948 61946 38976 68750
rect 39040 68338 39068 69158
rect 39028 68332 39080 68338
rect 39028 68274 39080 68280
rect 39316 68270 39344 71200
rect 41420 69216 41472 69222
rect 41420 69158 41472 69164
rect 41432 68882 41460 69158
rect 41892 68882 41920 71200
rect 42892 69216 42944 69222
rect 42892 69158 42944 69164
rect 42904 68882 42932 69158
rect 43180 68882 43208 71200
rect 41420 68876 41472 68882
rect 41420 68818 41472 68824
rect 41880 68876 41932 68882
rect 41880 68818 41932 68824
rect 42892 68876 42944 68882
rect 42892 68818 42944 68824
rect 43168 68876 43220 68882
rect 43168 68818 43220 68824
rect 39856 68808 39908 68814
rect 39856 68750 39908 68756
rect 39764 68672 39816 68678
rect 39764 68614 39816 68620
rect 39776 68406 39804 68614
rect 39868 68406 39896 68750
rect 41420 68740 41472 68746
rect 41420 68682 41472 68688
rect 42800 68740 42852 68746
rect 42800 68682 42852 68688
rect 39764 68400 39816 68406
rect 39764 68342 39816 68348
rect 39856 68400 39908 68406
rect 39856 68342 39908 68348
rect 39304 68264 39356 68270
rect 39304 68206 39356 68212
rect 41432 67930 41460 68682
rect 42616 68672 42668 68678
rect 42616 68614 42668 68620
rect 42628 68474 42656 68614
rect 42812 68474 42840 68682
rect 42616 68468 42668 68474
rect 42616 68410 42668 68416
rect 42800 68468 42852 68474
rect 42800 68410 42852 68416
rect 42708 68196 42760 68202
rect 42708 68138 42760 68144
rect 41420 67924 41472 67930
rect 41420 67866 41472 67872
rect 41328 67720 41380 67726
rect 41328 67662 41380 67668
rect 41340 67182 41368 67662
rect 40960 67176 41012 67182
rect 40960 67118 41012 67124
rect 41328 67176 41380 67182
rect 41328 67118 41380 67124
rect 38936 61940 38988 61946
rect 38936 61882 38988 61888
rect 39948 61192 40000 61198
rect 39948 61134 40000 61140
rect 38752 61124 38804 61130
rect 38752 61066 38804 61072
rect 38660 60716 38712 60722
rect 38660 60658 38712 60664
rect 38672 60314 38700 60658
rect 38660 60308 38712 60314
rect 38660 60250 38712 60256
rect 38764 58614 38792 61066
rect 39856 60716 39908 60722
rect 39856 60658 39908 60664
rect 39212 60512 39264 60518
rect 39212 60454 39264 60460
rect 38844 60172 38896 60178
rect 38844 60114 38896 60120
rect 38856 59022 38884 60114
rect 38936 60104 38988 60110
rect 38936 60046 38988 60052
rect 38844 59016 38896 59022
rect 38844 58958 38896 58964
rect 38856 58886 38884 58958
rect 38844 58880 38896 58886
rect 38844 58822 38896 58828
rect 38752 58608 38804 58614
rect 38752 58550 38804 58556
rect 38660 58336 38712 58342
rect 38660 58278 38712 58284
rect 38672 57934 38700 58278
rect 38660 57928 38712 57934
rect 38660 57870 38712 57876
rect 38672 57390 38700 57870
rect 38764 57526 38792 58550
rect 38856 58290 38884 58822
rect 38948 58410 38976 60046
rect 39224 59566 39252 60454
rect 39672 60104 39724 60110
rect 39672 60046 39724 60052
rect 39684 59634 39712 60046
rect 39672 59628 39724 59634
rect 39672 59570 39724 59576
rect 39212 59560 39264 59566
rect 39212 59502 39264 59508
rect 39120 59424 39172 59430
rect 39120 59366 39172 59372
rect 39132 59090 39160 59366
rect 39120 59084 39172 59090
rect 39120 59026 39172 59032
rect 39132 58614 39160 59026
rect 39120 58608 39172 58614
rect 39120 58550 39172 58556
rect 39224 58546 39252 59502
rect 39684 59090 39712 59570
rect 39868 59226 39896 60658
rect 39960 60178 39988 61134
rect 40132 61124 40184 61130
rect 40132 61066 40184 61072
rect 40144 60858 40172 61066
rect 40132 60852 40184 60858
rect 40132 60794 40184 60800
rect 40132 60716 40184 60722
rect 40132 60658 40184 60664
rect 40144 60314 40172 60658
rect 40132 60308 40184 60314
rect 40132 60250 40184 60256
rect 39948 60172 40000 60178
rect 39948 60114 40000 60120
rect 40132 60104 40184 60110
rect 39960 60052 40132 60058
rect 39960 60046 40184 60052
rect 39960 60030 40172 60046
rect 40224 60036 40276 60042
rect 39856 59220 39908 59226
rect 39856 59162 39908 59168
rect 39672 59084 39724 59090
rect 39672 59026 39724 59032
rect 39684 58682 39712 59026
rect 39960 59022 39988 60030
rect 40224 59978 40276 59984
rect 40236 59090 40264 59978
rect 40224 59084 40276 59090
rect 40224 59026 40276 59032
rect 39948 59016 40000 59022
rect 39948 58958 40000 58964
rect 39960 58886 39988 58958
rect 40236 58954 40264 59026
rect 40316 59016 40368 59022
rect 40316 58958 40368 58964
rect 40776 59016 40828 59022
rect 40776 58958 40828 58964
rect 40224 58948 40276 58954
rect 40224 58890 40276 58896
rect 39948 58880 40000 58886
rect 39948 58822 40000 58828
rect 39672 58676 39724 58682
rect 39672 58618 39724 58624
rect 39960 58546 39988 58822
rect 39212 58540 39264 58546
rect 39212 58482 39264 58488
rect 39948 58540 40000 58546
rect 39948 58482 40000 58488
rect 40236 58478 40264 58890
rect 40328 58546 40356 58958
rect 40316 58540 40368 58546
rect 40316 58482 40368 58488
rect 40224 58472 40276 58478
rect 40224 58414 40276 58420
rect 38936 58404 38988 58410
rect 38936 58346 38988 58352
rect 38856 58262 38976 58290
rect 38844 57928 38896 57934
rect 38844 57870 38896 57876
rect 38752 57520 38804 57526
rect 38752 57462 38804 57468
rect 38856 57458 38884 57870
rect 38844 57452 38896 57458
rect 38844 57394 38896 57400
rect 38660 57384 38712 57390
rect 38948 57338 38976 58262
rect 39028 58064 39080 58070
rect 39028 58006 39080 58012
rect 38660 57326 38712 57332
rect 38856 57310 38976 57338
rect 38856 57050 38884 57310
rect 38936 57248 38988 57254
rect 38936 57190 38988 57196
rect 38844 57044 38896 57050
rect 38844 56986 38896 56992
rect 38948 56846 38976 57190
rect 38936 56840 38988 56846
rect 38936 56782 38988 56788
rect 38752 56704 38804 56710
rect 38752 56646 38804 56652
rect 38844 56704 38896 56710
rect 38844 56646 38896 56652
rect 38764 56370 38792 56646
rect 38752 56364 38804 56370
rect 38752 56306 38804 56312
rect 38764 55826 38792 56306
rect 38856 56302 38884 56646
rect 38844 56296 38896 56302
rect 39040 56250 39068 58006
rect 40788 57594 40816 58958
rect 40776 57588 40828 57594
rect 40776 57530 40828 57536
rect 39120 57384 39172 57390
rect 39120 57326 39172 57332
rect 38844 56238 38896 56244
rect 38948 56222 39068 56250
rect 38752 55820 38804 55826
rect 38752 55762 38804 55768
rect 38948 55758 38976 56222
rect 39132 56114 39160 57326
rect 40788 56914 40816 57530
rect 40776 56908 40828 56914
rect 40776 56850 40828 56856
rect 40500 56704 40552 56710
rect 40500 56646 40552 56652
rect 40512 56370 40540 56646
rect 40684 56500 40736 56506
rect 40684 56442 40736 56448
rect 40696 56370 40724 56442
rect 40500 56364 40552 56370
rect 40500 56306 40552 56312
rect 40684 56364 40736 56370
rect 40684 56306 40736 56312
rect 39040 56086 39160 56114
rect 39040 55758 39068 56086
rect 39120 55820 39172 55826
rect 39120 55762 39172 55768
rect 38936 55752 38988 55758
rect 38936 55694 38988 55700
rect 39028 55752 39080 55758
rect 39028 55694 39080 55700
rect 38660 55616 38712 55622
rect 38660 55558 38712 55564
rect 38672 54874 38700 55558
rect 38948 55298 38976 55694
rect 39040 55418 39068 55694
rect 39028 55412 39080 55418
rect 39028 55354 39080 55360
rect 38948 55270 39068 55298
rect 39132 55282 39160 55762
rect 40788 55758 40816 56850
rect 40776 55752 40828 55758
rect 40776 55694 40828 55700
rect 40500 55684 40552 55690
rect 40500 55626 40552 55632
rect 40512 55418 40540 55626
rect 40500 55412 40552 55418
rect 40500 55354 40552 55360
rect 39040 55214 39068 55270
rect 39120 55276 39172 55282
rect 39120 55218 39172 55224
rect 39028 55208 39080 55214
rect 39028 55150 39080 55156
rect 38660 54868 38712 54874
rect 38660 54810 38712 54816
rect 38936 54664 38988 54670
rect 38936 54606 38988 54612
rect 38948 53990 38976 54606
rect 40040 54188 40092 54194
rect 40040 54130 40092 54136
rect 38936 53984 38988 53990
rect 38936 53926 38988 53932
rect 38844 53508 38896 53514
rect 38844 53450 38896 53456
rect 38856 51406 38884 53450
rect 38660 51400 38712 51406
rect 38660 51342 38712 51348
rect 38844 51400 38896 51406
rect 38844 51342 38896 51348
rect 38568 50312 38620 50318
rect 38568 50254 38620 50260
rect 38292 49904 38344 49910
rect 38292 49846 38344 49852
rect 38304 49230 38332 49846
rect 38292 49224 38344 49230
rect 38292 49166 38344 49172
rect 38120 48286 38240 48314
rect 37924 48068 37976 48074
rect 37924 48010 37976 48016
rect 38016 48068 38068 48074
rect 38016 48010 38068 48016
rect 37832 47660 37884 47666
rect 37832 47602 37884 47608
rect 37844 47190 37872 47602
rect 37832 47184 37884 47190
rect 37832 47126 37884 47132
rect 37936 46986 37964 48010
rect 38028 47258 38056 48010
rect 38016 47252 38068 47258
rect 38016 47194 38068 47200
rect 38016 47048 38068 47054
rect 38016 46990 38068 46996
rect 38108 47048 38160 47054
rect 38108 46990 38160 46996
rect 37924 46980 37976 46986
rect 37924 46922 37976 46928
rect 37740 45824 37792 45830
rect 37740 45766 37792 45772
rect 37648 42628 37700 42634
rect 37648 42570 37700 42576
rect 37648 42016 37700 42022
rect 37648 41958 37700 41964
rect 37660 41857 37688 41958
rect 37646 41848 37702 41857
rect 37646 41783 37702 41792
rect 37752 41562 37780 45766
rect 37936 43790 37964 46922
rect 38028 45286 38056 46990
rect 38016 45280 38068 45286
rect 38016 45222 38068 45228
rect 38028 44946 38056 45222
rect 38016 44940 38068 44946
rect 38016 44882 38068 44888
rect 38120 43790 38148 46990
rect 38212 46934 38240 48286
rect 38212 46906 38332 46934
rect 38200 46504 38252 46510
rect 38200 46446 38252 46452
rect 37924 43784 37976 43790
rect 37924 43726 37976 43732
rect 38108 43784 38160 43790
rect 38108 43726 38160 43732
rect 37832 43308 37884 43314
rect 37832 43250 37884 43256
rect 37844 42566 37872 43250
rect 37936 42702 37964 43726
rect 37924 42696 37976 42702
rect 37924 42638 37976 42644
rect 38016 42628 38068 42634
rect 38016 42570 38068 42576
rect 37832 42560 37884 42566
rect 37832 42502 37884 42508
rect 37568 41534 37780 41562
rect 37464 41472 37516 41478
rect 37464 41414 37516 41420
rect 37568 41206 37596 41534
rect 37740 41472 37792 41478
rect 37646 41440 37702 41449
rect 37740 41414 37792 41420
rect 37646 41375 37702 41384
rect 37556 41200 37608 41206
rect 37556 41142 37608 41148
rect 37464 41132 37516 41138
rect 37464 41074 37516 41080
rect 37372 40520 37424 40526
rect 37372 40462 37424 40468
rect 37384 38418 37412 40462
rect 37372 38412 37424 38418
rect 37372 38354 37424 38360
rect 37476 37942 37504 41074
rect 37660 41018 37688 41375
rect 37752 41138 37780 41414
rect 37844 41138 37872 42502
rect 37924 42288 37976 42294
rect 37924 42230 37976 42236
rect 37740 41132 37792 41138
rect 37740 41074 37792 41080
rect 37832 41132 37884 41138
rect 37832 41074 37884 41080
rect 37556 40996 37608 41002
rect 37660 40990 37872 41018
rect 37556 40938 37608 40944
rect 37568 40662 37596 40938
rect 37648 40928 37700 40934
rect 37648 40870 37700 40876
rect 37660 40662 37688 40870
rect 37844 40730 37872 40990
rect 37832 40724 37884 40730
rect 37832 40666 37884 40672
rect 37556 40656 37608 40662
rect 37556 40598 37608 40604
rect 37648 40656 37700 40662
rect 37648 40598 37700 40604
rect 37740 40452 37792 40458
rect 37740 40394 37792 40400
rect 37648 39840 37700 39846
rect 37648 39782 37700 39788
rect 37660 39574 37688 39782
rect 37648 39568 37700 39574
rect 37648 39510 37700 39516
rect 37648 38344 37700 38350
rect 37648 38286 37700 38292
rect 37464 37936 37516 37942
rect 37464 37878 37516 37884
rect 37372 36780 37424 36786
rect 37372 36722 37424 36728
rect 37280 35692 37332 35698
rect 37280 35634 37332 35640
rect 37188 34468 37240 34474
rect 37188 34410 37240 34416
rect 37292 33998 37320 35634
rect 37384 35290 37412 36722
rect 37372 35284 37424 35290
rect 37372 35226 37424 35232
rect 37476 35018 37504 37878
rect 37556 37868 37608 37874
rect 37556 37810 37608 37816
rect 37568 37466 37596 37810
rect 37556 37460 37608 37466
rect 37556 37402 37608 37408
rect 37464 35012 37516 35018
rect 37464 34954 37516 34960
rect 37280 33992 37332 33998
rect 37280 33934 37332 33940
rect 37004 33040 37056 33046
rect 37004 32982 37056 32988
rect 37292 32978 37320 33934
rect 37372 33380 37424 33386
rect 37372 33322 37424 33328
rect 37280 32972 37332 32978
rect 37280 32914 37332 32920
rect 37384 32910 37412 33322
rect 37476 32910 37504 34954
rect 37372 32904 37424 32910
rect 37372 32846 37424 32852
rect 37464 32904 37516 32910
rect 37464 32846 37516 32852
rect 37660 32502 37688 38286
rect 37752 34678 37780 40394
rect 37844 40050 37872 40666
rect 37832 40044 37884 40050
rect 37832 39986 37884 39992
rect 37844 39438 37872 39986
rect 37936 39914 37964 42230
rect 38028 41414 38056 42570
rect 38106 41576 38162 41585
rect 38106 41511 38108 41520
rect 38160 41511 38162 41520
rect 38108 41482 38160 41488
rect 38028 41386 38148 41414
rect 38120 41290 38148 41386
rect 38028 41262 38148 41290
rect 38028 40390 38056 41262
rect 38108 41132 38160 41138
rect 38108 41074 38160 41080
rect 38016 40384 38068 40390
rect 38016 40326 38068 40332
rect 37924 39908 37976 39914
rect 37924 39850 37976 39856
rect 37832 39432 37884 39438
rect 37832 39374 37884 39380
rect 37844 36922 37872 39374
rect 37832 36916 37884 36922
rect 37832 36858 37884 36864
rect 37924 36168 37976 36174
rect 37924 36110 37976 36116
rect 37936 35834 37964 36110
rect 37924 35828 37976 35834
rect 37924 35770 37976 35776
rect 38028 35698 38056 40326
rect 38120 40186 38148 41074
rect 38108 40180 38160 40186
rect 38108 40122 38160 40128
rect 38212 40118 38240 46446
rect 38304 46442 38332 46906
rect 38568 46572 38620 46578
rect 38568 46514 38620 46520
rect 38292 46436 38344 46442
rect 38292 46378 38344 46384
rect 38476 43648 38528 43654
rect 38476 43590 38528 43596
rect 38384 41676 38436 41682
rect 38384 41618 38436 41624
rect 38292 41608 38344 41614
rect 38292 41550 38344 41556
rect 38304 40916 38332 41550
rect 38396 41138 38424 41618
rect 38384 41132 38436 41138
rect 38384 41074 38436 41080
rect 38384 40928 38436 40934
rect 38304 40888 38384 40916
rect 38384 40870 38436 40876
rect 38488 40594 38516 43590
rect 38476 40588 38528 40594
rect 38476 40530 38528 40536
rect 38200 40112 38252 40118
rect 38200 40054 38252 40060
rect 38384 39908 38436 39914
rect 38384 39850 38436 39856
rect 38200 39296 38252 39302
rect 38200 39238 38252 39244
rect 38212 38962 38240 39238
rect 38200 38956 38252 38962
rect 38200 38898 38252 38904
rect 38396 38350 38424 39850
rect 38476 39432 38528 39438
rect 38476 39374 38528 39380
rect 38488 39098 38516 39374
rect 38476 39092 38528 39098
rect 38476 39034 38528 39040
rect 38384 38344 38436 38350
rect 38384 38286 38436 38292
rect 38384 36916 38436 36922
rect 38384 36858 38436 36864
rect 38396 36786 38424 36858
rect 38384 36780 38436 36786
rect 38384 36722 38436 36728
rect 38016 35692 38068 35698
rect 38016 35634 38068 35640
rect 38016 34944 38068 34950
rect 38016 34886 38068 34892
rect 38108 34944 38160 34950
rect 38108 34886 38160 34892
rect 37740 34672 37792 34678
rect 37740 34614 37792 34620
rect 38028 34610 38056 34886
rect 38016 34604 38068 34610
rect 38016 34546 38068 34552
rect 37832 34400 37884 34406
rect 37832 34342 37884 34348
rect 37372 32496 37424 32502
rect 37372 32438 37424 32444
rect 37648 32496 37700 32502
rect 37648 32438 37700 32444
rect 37384 31822 37412 32438
rect 37372 31816 37424 31822
rect 37372 31758 37424 31764
rect 37384 30326 37412 31758
rect 37844 31754 37872 34342
rect 38120 33998 38148 34886
rect 38108 33992 38160 33998
rect 38108 33934 38160 33940
rect 38384 32768 38436 32774
rect 38384 32710 38436 32716
rect 38396 32434 38424 32710
rect 38384 32428 38436 32434
rect 38384 32370 38436 32376
rect 38292 32360 38344 32366
rect 38292 32302 38344 32308
rect 38108 32224 38160 32230
rect 38108 32166 38160 32172
rect 37832 31748 37884 31754
rect 37832 31690 37884 31696
rect 37844 31346 37872 31690
rect 37832 31340 37884 31346
rect 37832 31282 37884 31288
rect 37556 31136 37608 31142
rect 37556 31078 37608 31084
rect 37568 30802 37596 31078
rect 37556 30796 37608 30802
rect 37556 30738 37608 30744
rect 37372 30320 37424 30326
rect 37372 30262 37424 30268
rect 37384 29646 37412 30262
rect 37372 29640 37424 29646
rect 37372 29582 37424 29588
rect 38120 29238 38148 32166
rect 38304 32026 38332 32302
rect 38292 32020 38344 32026
rect 38292 31962 38344 31968
rect 38200 30660 38252 30666
rect 38200 30602 38252 30608
rect 38212 30394 38240 30602
rect 38200 30388 38252 30394
rect 38200 30330 38252 30336
rect 38384 30252 38436 30258
rect 38384 30194 38436 30200
rect 38396 29850 38424 30194
rect 38384 29844 38436 29850
rect 38384 29786 38436 29792
rect 38108 29232 38160 29238
rect 38108 29174 38160 29180
rect 38200 29164 38252 29170
rect 38200 29106 38252 29112
rect 37924 28960 37976 28966
rect 37924 28902 37976 28908
rect 37936 28490 37964 28902
rect 37924 28484 37976 28490
rect 37924 28426 37976 28432
rect 38212 28422 38240 29106
rect 38200 28416 38252 28422
rect 38200 28358 38252 28364
rect 38488 27606 38516 39034
rect 38580 38010 38608 46514
rect 38672 46374 38700 51342
rect 38752 51264 38804 51270
rect 38752 51206 38804 51212
rect 38764 50794 38792 51206
rect 38752 50788 38804 50794
rect 38752 50730 38804 50736
rect 38752 47456 38804 47462
rect 38752 47398 38804 47404
rect 38660 46368 38712 46374
rect 38660 46310 38712 46316
rect 38660 43852 38712 43858
rect 38660 43794 38712 43800
rect 38672 43722 38700 43794
rect 38660 43716 38712 43722
rect 38660 43658 38712 43664
rect 38672 43382 38700 43658
rect 38660 43376 38712 43382
rect 38660 43318 38712 43324
rect 38660 41608 38712 41614
rect 38660 41550 38712 41556
rect 38672 41177 38700 41550
rect 38658 41168 38714 41177
rect 38658 41103 38714 41112
rect 38660 41064 38712 41070
rect 38660 41006 38712 41012
rect 38672 40458 38700 41006
rect 38764 40474 38792 47398
rect 38856 43858 38884 51342
rect 38948 47054 38976 53926
rect 39396 53576 39448 53582
rect 39396 53518 39448 53524
rect 39408 51074 39436 53518
rect 39488 53440 39540 53446
rect 39488 53382 39540 53388
rect 39500 53106 39528 53382
rect 40052 53242 40080 54130
rect 40776 53984 40828 53990
rect 40776 53926 40828 53932
rect 40224 53508 40276 53514
rect 40224 53450 40276 53456
rect 40040 53236 40092 53242
rect 40040 53178 40092 53184
rect 39488 53100 39540 53106
rect 39488 53042 39540 53048
rect 40236 51074 40264 53450
rect 40788 53174 40816 53926
rect 40776 53168 40828 53174
rect 40776 53110 40828 53116
rect 39408 51046 39528 51074
rect 40236 51046 40448 51074
rect 39500 50930 39528 51046
rect 39488 50924 39540 50930
rect 39488 50866 39540 50872
rect 39500 48278 39528 50866
rect 39672 50312 39724 50318
rect 39672 50254 39724 50260
rect 39684 49842 39712 50254
rect 39672 49836 39724 49842
rect 39672 49778 39724 49784
rect 39684 49230 39712 49778
rect 40040 49428 40092 49434
rect 40040 49370 40092 49376
rect 39672 49224 39724 49230
rect 39672 49166 39724 49172
rect 39488 48272 39540 48278
rect 39488 48214 39540 48220
rect 39396 47660 39448 47666
rect 39396 47602 39448 47608
rect 39408 47258 39436 47602
rect 39684 47598 39712 49166
rect 40052 48142 40080 49370
rect 40132 49360 40184 49366
rect 40132 49302 40184 49308
rect 40144 48210 40172 49302
rect 40224 49088 40276 49094
rect 40224 49030 40276 49036
rect 40316 49088 40368 49094
rect 40316 49030 40368 49036
rect 40236 48686 40264 49030
rect 40224 48680 40276 48686
rect 40224 48622 40276 48628
rect 40132 48204 40184 48210
rect 40132 48146 40184 48152
rect 40040 48136 40092 48142
rect 40040 48078 40092 48084
rect 40224 48136 40276 48142
rect 40224 48078 40276 48084
rect 39856 48000 39908 48006
rect 39856 47942 39908 47948
rect 39672 47592 39724 47598
rect 39672 47534 39724 47540
rect 39396 47252 39448 47258
rect 39396 47194 39448 47200
rect 38936 47048 38988 47054
rect 38936 46990 38988 46996
rect 39028 46436 39080 46442
rect 39028 46378 39080 46384
rect 38844 43852 38896 43858
rect 38844 43794 38896 43800
rect 38936 43784 38988 43790
rect 38936 43726 38988 43732
rect 38844 43716 38896 43722
rect 38844 43658 38896 43664
rect 38856 43450 38884 43658
rect 38844 43444 38896 43450
rect 38844 43386 38896 43392
rect 38844 43240 38896 43246
rect 38844 43182 38896 43188
rect 38856 42906 38884 43182
rect 38844 42900 38896 42906
rect 38844 42842 38896 42848
rect 38948 42090 38976 43726
rect 39040 42158 39068 46378
rect 39120 46368 39172 46374
rect 39120 46310 39172 46316
rect 39028 42152 39080 42158
rect 39028 42094 39080 42100
rect 38936 42084 38988 42090
rect 38936 42026 38988 42032
rect 38844 42016 38896 42022
rect 38844 41958 38896 41964
rect 38856 41614 38884 41958
rect 39028 41744 39080 41750
rect 39026 41712 39028 41721
rect 39080 41712 39082 41721
rect 39026 41647 39082 41656
rect 38844 41608 38896 41614
rect 38844 41550 38896 41556
rect 38936 41540 38988 41546
rect 38936 41482 38988 41488
rect 38948 41002 38976 41482
rect 39028 41472 39080 41478
rect 39028 41414 39080 41420
rect 39040 41206 39068 41414
rect 39028 41200 39080 41206
rect 39028 41142 39080 41148
rect 38936 40996 38988 41002
rect 38936 40938 38988 40944
rect 39028 40588 39080 40594
rect 39028 40530 39080 40536
rect 38660 40452 38712 40458
rect 38764 40446 38884 40474
rect 38660 40394 38712 40400
rect 38752 40384 38804 40390
rect 38752 40326 38804 40332
rect 38764 39438 38792 40326
rect 38856 39506 38884 40446
rect 39040 39828 39068 40530
rect 39132 40526 39160 46310
rect 39868 45558 39896 47942
rect 39948 47660 40000 47666
rect 39948 47602 40000 47608
rect 39960 46986 39988 47602
rect 40040 47456 40092 47462
rect 40040 47398 40092 47404
rect 40052 47138 40080 47398
rect 40236 47258 40264 48078
rect 40224 47252 40276 47258
rect 40224 47194 40276 47200
rect 40052 47122 40172 47138
rect 40052 47116 40184 47122
rect 40052 47110 40132 47116
rect 40052 46986 40080 47110
rect 40132 47058 40184 47064
rect 39948 46980 40000 46986
rect 39948 46922 40000 46928
rect 40040 46980 40092 46986
rect 40040 46922 40092 46928
rect 40236 46646 40264 47194
rect 40224 46640 40276 46646
rect 40224 46582 40276 46588
rect 39948 46504 40000 46510
rect 39948 46446 40000 46452
rect 39856 45552 39908 45558
rect 39856 45494 39908 45500
rect 39856 43444 39908 43450
rect 39856 43386 39908 43392
rect 39396 43308 39448 43314
rect 39396 43250 39448 43256
rect 39408 42090 39436 43250
rect 39868 42770 39896 43386
rect 39960 42906 39988 46446
rect 40132 46368 40184 46374
rect 40132 46310 40184 46316
rect 40144 45966 40172 46310
rect 40040 45960 40092 45966
rect 40040 45902 40092 45908
rect 40132 45960 40184 45966
rect 40132 45902 40184 45908
rect 40052 45082 40080 45902
rect 40040 45076 40092 45082
rect 40040 45018 40092 45024
rect 39948 42900 40000 42906
rect 39948 42842 40000 42848
rect 39856 42764 39908 42770
rect 39856 42706 39908 42712
rect 39764 42560 39816 42566
rect 39764 42502 39816 42508
rect 39776 42226 39804 42502
rect 39580 42220 39632 42226
rect 39580 42162 39632 42168
rect 39764 42220 39816 42226
rect 39764 42162 39816 42168
rect 39212 42084 39264 42090
rect 39212 42026 39264 42032
rect 39396 42084 39448 42090
rect 39396 42026 39448 42032
rect 39120 40520 39172 40526
rect 39120 40462 39172 40468
rect 39224 40118 39252 42026
rect 39592 41682 39620 42162
rect 39580 41676 39632 41682
rect 39580 41618 39632 41624
rect 39960 41414 39988 42842
rect 40328 42702 40356 49030
rect 40420 43994 40448 51046
rect 40500 50516 40552 50522
rect 40500 50458 40552 50464
rect 40408 43988 40460 43994
rect 40408 43930 40460 43936
rect 40512 43790 40540 50458
rect 40972 48634 41000 67118
rect 41236 61056 41288 61062
rect 41236 60998 41288 61004
rect 41248 60042 41276 60998
rect 42720 60110 42748 68138
rect 44468 64874 44496 71200
rect 45192 69216 45244 69222
rect 45192 69158 45244 69164
rect 45204 68338 45232 69158
rect 45376 68672 45428 68678
rect 45376 68614 45428 68620
rect 45388 68406 45416 68614
rect 45376 68400 45428 68406
rect 45376 68342 45428 68348
rect 45192 68332 45244 68338
rect 45192 68274 45244 68280
rect 45756 68270 45784 71200
rect 46480 69420 46532 69426
rect 46480 69362 46532 69368
rect 46112 69216 46164 69222
rect 46112 69158 46164 69164
rect 46124 68882 46152 69158
rect 46112 68876 46164 68882
rect 46112 68818 46164 68824
rect 45744 68264 45796 68270
rect 45744 68206 45796 68212
rect 46492 66026 46520 69362
rect 46572 69216 46624 69222
rect 46572 69158 46624 69164
rect 46584 68882 46612 69158
rect 47044 68882 47072 71200
rect 46572 68876 46624 68882
rect 46572 68818 46624 68824
rect 47032 68876 47084 68882
rect 47032 68818 47084 68824
rect 46480 66020 46532 66026
rect 46480 65962 46532 65968
rect 44192 64846 44496 64874
rect 44192 62966 44220 64846
rect 44180 62960 44232 62966
rect 44180 62902 44232 62908
rect 42708 60104 42760 60110
rect 42708 60046 42760 60052
rect 41236 60036 41288 60042
rect 41236 59978 41288 59984
rect 44088 60036 44140 60042
rect 44088 59978 44140 59984
rect 42984 59968 43036 59974
rect 42984 59910 43036 59916
rect 42996 59634 43024 59910
rect 44100 59770 44128 59978
rect 44088 59764 44140 59770
rect 44088 59706 44140 59712
rect 41604 59628 41656 59634
rect 41604 59570 41656 59576
rect 41696 59628 41748 59634
rect 41696 59570 41748 59576
rect 42984 59628 43036 59634
rect 42984 59570 43036 59576
rect 43536 59628 43588 59634
rect 43536 59570 43588 59576
rect 44180 59628 44232 59634
rect 44180 59570 44232 59576
rect 41512 59560 41564 59566
rect 41512 59502 41564 59508
rect 41420 59424 41472 59430
rect 41420 59366 41472 59372
rect 41236 58948 41288 58954
rect 41236 58890 41288 58896
rect 41248 58682 41276 58890
rect 41236 58676 41288 58682
rect 41236 58618 41288 58624
rect 41432 58546 41460 59366
rect 41524 58614 41552 59502
rect 41616 59226 41644 59570
rect 41604 59220 41656 59226
rect 41604 59162 41656 59168
rect 41512 58608 41564 58614
rect 41512 58550 41564 58556
rect 41420 58540 41472 58546
rect 41420 58482 41472 58488
rect 41524 58426 41552 58550
rect 41616 58546 41644 59162
rect 41604 58540 41656 58546
rect 41604 58482 41656 58488
rect 41708 58426 41736 59570
rect 42616 59560 42668 59566
rect 42616 59502 42668 59508
rect 42628 59090 42656 59502
rect 42708 59492 42760 59498
rect 42708 59434 42760 59440
rect 42616 59084 42668 59090
rect 42616 59026 42668 59032
rect 42720 59022 42748 59434
rect 42708 59016 42760 59022
rect 42708 58958 42760 58964
rect 41432 58398 41552 58426
rect 41616 58398 41736 58426
rect 42720 58410 42748 58958
rect 42996 58954 43024 59570
rect 43548 59514 43576 59570
rect 43088 59486 43576 59514
rect 43088 59430 43116 59486
rect 43076 59424 43128 59430
rect 43076 59366 43128 59372
rect 43168 59424 43220 59430
rect 43168 59366 43220 59372
rect 42984 58948 43036 58954
rect 42984 58890 43036 58896
rect 42996 58546 43024 58890
rect 42984 58540 43036 58546
rect 42984 58482 43036 58488
rect 43180 58478 43208 59366
rect 44192 59226 44220 59570
rect 44180 59220 44232 59226
rect 44180 59162 44232 59168
rect 43444 59016 43496 59022
rect 43444 58958 43496 58964
rect 43456 58478 43484 58958
rect 43168 58472 43220 58478
rect 43168 58414 43220 58420
rect 43444 58472 43496 58478
rect 43444 58414 43496 58420
rect 43720 58472 43772 58478
rect 43720 58414 43772 58420
rect 43904 58472 43956 58478
rect 43904 58414 43956 58420
rect 42708 58404 42760 58410
rect 41432 58342 41460 58398
rect 41616 58342 41644 58398
rect 42708 58346 42760 58352
rect 41420 58336 41472 58342
rect 41420 58278 41472 58284
rect 41604 58336 41656 58342
rect 41604 58278 41656 58284
rect 41328 57452 41380 57458
rect 41328 57394 41380 57400
rect 41144 57248 41196 57254
rect 41144 57190 41196 57196
rect 41156 56778 41184 57190
rect 41144 56772 41196 56778
rect 41144 56714 41196 56720
rect 41340 56506 41368 57394
rect 41328 56500 41380 56506
rect 41328 56442 41380 56448
rect 41328 55276 41380 55282
rect 41328 55218 41380 55224
rect 41340 54738 41368 55218
rect 41328 54732 41380 54738
rect 41328 54674 41380 54680
rect 41340 54058 41368 54674
rect 41432 54602 41460 58278
rect 41616 56234 41644 58278
rect 43076 57860 43128 57866
rect 43076 57802 43128 57808
rect 42984 57452 43036 57458
rect 42984 57394 43036 57400
rect 42800 57384 42852 57390
rect 42800 57326 42852 57332
rect 42892 57384 42944 57390
rect 42892 57326 42944 57332
rect 42616 57248 42668 57254
rect 42616 57190 42668 57196
rect 42524 56840 42576 56846
rect 42524 56782 42576 56788
rect 42156 56704 42208 56710
rect 42156 56646 42208 56652
rect 42168 56302 42196 56646
rect 42156 56296 42208 56302
rect 42156 56238 42208 56244
rect 41604 56228 41656 56234
rect 41604 56170 41656 56176
rect 42432 56160 42484 56166
rect 42432 56102 42484 56108
rect 42444 55214 42472 56102
rect 42536 55282 42564 56782
rect 42628 56234 42656 57190
rect 42812 56302 42840 57326
rect 42904 57050 42932 57326
rect 42892 57044 42944 57050
rect 42892 56986 42944 56992
rect 42904 56438 42932 56986
rect 42892 56432 42944 56438
rect 42892 56374 42944 56380
rect 42800 56296 42852 56302
rect 42800 56238 42852 56244
rect 42616 56228 42668 56234
rect 42616 56170 42668 56176
rect 42996 56166 43024 57394
rect 43088 56914 43116 57802
rect 43076 56908 43128 56914
rect 43076 56850 43128 56856
rect 43180 56794 43208 58414
rect 43732 57458 43760 58414
rect 43916 58138 43944 58414
rect 44272 58336 44324 58342
rect 44272 58278 44324 58284
rect 43904 58132 43956 58138
rect 43904 58074 43956 58080
rect 44284 57934 44312 58278
rect 44272 57928 44324 57934
rect 44272 57870 44324 57876
rect 46388 57792 46440 57798
rect 46388 57734 46440 57740
rect 46400 57458 46428 57734
rect 43720 57452 43772 57458
rect 43720 57394 43772 57400
rect 46388 57452 46440 57458
rect 46388 57394 46440 57400
rect 43088 56766 43208 56794
rect 45376 56840 45428 56846
rect 45376 56782 45428 56788
rect 46848 56840 46900 56846
rect 46848 56782 46900 56788
rect 43352 56772 43404 56778
rect 42984 56160 43036 56166
rect 42984 56102 43036 56108
rect 42524 55276 42576 55282
rect 42524 55218 42576 55224
rect 42432 55208 42484 55214
rect 42432 55150 42484 55156
rect 43088 54670 43116 56766
rect 43352 56714 43404 56720
rect 43364 56506 43392 56714
rect 45192 56704 45244 56710
rect 45192 56646 45244 56652
rect 43352 56500 43404 56506
rect 43352 56442 43404 56448
rect 45204 56370 45232 56646
rect 43536 56364 43588 56370
rect 43536 56306 43588 56312
rect 45192 56364 45244 56370
rect 45192 56306 45244 56312
rect 43168 55276 43220 55282
rect 43168 55218 43220 55224
rect 43076 54664 43128 54670
rect 43076 54606 43128 54612
rect 41420 54596 41472 54602
rect 41420 54538 41472 54544
rect 41604 54596 41656 54602
rect 41604 54538 41656 54544
rect 41420 54188 41472 54194
rect 41420 54130 41472 54136
rect 41328 54052 41380 54058
rect 41328 53994 41380 54000
rect 41236 53236 41288 53242
rect 41236 53178 41288 53184
rect 41248 52018 41276 53178
rect 41236 52012 41288 52018
rect 41236 51954 41288 51960
rect 41248 51814 41276 51954
rect 41236 51808 41288 51814
rect 41236 51750 41288 51756
rect 41052 50924 41104 50930
rect 41052 50866 41104 50872
rect 41064 50522 41092 50866
rect 41052 50516 41104 50522
rect 41052 50458 41104 50464
rect 41340 50318 41368 53994
rect 41432 53582 41460 54130
rect 41512 53984 41564 53990
rect 41512 53926 41564 53932
rect 41524 53650 41552 53926
rect 41512 53644 41564 53650
rect 41512 53586 41564 53592
rect 41420 53576 41472 53582
rect 41420 53518 41472 53524
rect 41616 53106 41644 54538
rect 41788 53508 41840 53514
rect 41788 53450 41840 53456
rect 41800 53242 41828 53450
rect 42892 53440 42944 53446
rect 42892 53382 42944 53388
rect 41788 53236 41840 53242
rect 41788 53178 41840 53184
rect 42800 53236 42852 53242
rect 42800 53178 42852 53184
rect 41604 53100 41656 53106
rect 41604 53042 41656 53048
rect 42616 53100 42668 53106
rect 42616 53042 42668 53048
rect 42708 53100 42760 53106
rect 42708 53042 42760 53048
rect 41420 53032 41472 53038
rect 41418 53000 41420 53009
rect 41472 53000 41474 53009
rect 41418 52935 41474 52944
rect 41604 52964 41656 52970
rect 41604 52906 41656 52912
rect 41616 52018 41644 52906
rect 42628 52562 42656 53042
rect 42720 53009 42748 53042
rect 42706 53000 42762 53009
rect 42706 52935 42762 52944
rect 42616 52556 42668 52562
rect 42616 52498 42668 52504
rect 42340 52420 42392 52426
rect 42340 52362 42392 52368
rect 41604 52012 41656 52018
rect 41604 51954 41656 51960
rect 41696 51944 41748 51950
rect 41696 51886 41748 51892
rect 41604 51876 41656 51882
rect 41604 51818 41656 51824
rect 41616 51542 41644 51818
rect 41708 51610 41736 51886
rect 41880 51876 41932 51882
rect 41880 51818 41932 51824
rect 41696 51604 41748 51610
rect 41696 51546 41748 51552
rect 41604 51536 41656 51542
rect 41892 51490 41920 51818
rect 41604 51478 41656 51484
rect 41800 51462 41920 51490
rect 41604 50788 41656 50794
rect 41604 50730 41656 50736
rect 41616 50386 41644 50730
rect 41800 50522 41828 51462
rect 42352 51406 42380 52362
rect 42812 52086 42840 53178
rect 42904 53174 42932 53382
rect 42892 53168 42944 53174
rect 42892 53110 42944 53116
rect 42892 52352 42944 52358
rect 42892 52294 42944 52300
rect 42800 52080 42852 52086
rect 42800 52022 42852 52028
rect 42812 51626 42840 52022
rect 42904 51814 42932 52294
rect 42892 51808 42944 51814
rect 42944 51768 43024 51796
rect 42892 51750 42944 51756
rect 42536 51598 42840 51626
rect 42536 51474 42564 51598
rect 42524 51468 42576 51474
rect 42524 51410 42576 51416
rect 42340 51400 42392 51406
rect 42340 51342 42392 51348
rect 42616 51400 42668 51406
rect 42616 51342 42668 51348
rect 41880 51332 41932 51338
rect 41880 51274 41932 51280
rect 41788 50516 41840 50522
rect 41788 50458 41840 50464
rect 41604 50380 41656 50386
rect 41604 50322 41656 50328
rect 41892 50318 41920 51274
rect 42628 50969 42656 51342
rect 42614 50960 42670 50969
rect 42614 50895 42670 50904
rect 42628 50794 42656 50895
rect 42812 50862 42840 51598
rect 42996 51406 43024 51768
rect 42984 51400 43036 51406
rect 42984 51342 43036 51348
rect 42800 50856 42852 50862
rect 42800 50798 42852 50804
rect 42616 50788 42668 50794
rect 42616 50730 42668 50736
rect 41328 50312 41380 50318
rect 41328 50254 41380 50260
rect 41880 50312 41932 50318
rect 41880 50254 41932 50260
rect 42432 50312 42484 50318
rect 42432 50254 42484 50260
rect 41340 49434 41368 50254
rect 41696 49904 41748 49910
rect 41696 49846 41748 49852
rect 41328 49428 41380 49434
rect 41328 49370 41380 49376
rect 41708 49366 41736 49846
rect 41696 49360 41748 49366
rect 41696 49302 41748 49308
rect 41420 49224 41472 49230
rect 41420 49166 41472 49172
rect 41696 49224 41748 49230
rect 41696 49166 41748 49172
rect 41432 48890 41460 49166
rect 41420 48884 41472 48890
rect 41420 48826 41472 48832
rect 41604 48748 41656 48754
rect 41604 48690 41656 48696
rect 41328 48680 41380 48686
rect 40972 48606 41092 48634
rect 41328 48622 41380 48628
rect 40684 48544 40736 48550
rect 40684 48486 40736 48492
rect 40960 48544 41012 48550
rect 40960 48486 41012 48492
rect 40696 48074 40724 48486
rect 40684 48068 40736 48074
rect 40684 48010 40736 48016
rect 40972 47666 41000 48486
rect 40960 47660 41012 47666
rect 40960 47602 41012 47608
rect 40972 47530 41000 47602
rect 40960 47524 41012 47530
rect 40960 47466 41012 47472
rect 40684 47456 40736 47462
rect 40684 47398 40736 47404
rect 40696 46578 40724 47398
rect 40972 47122 41000 47466
rect 40960 47116 41012 47122
rect 40960 47058 41012 47064
rect 40684 46572 40736 46578
rect 40684 46514 40736 46520
rect 41064 44470 41092 48606
rect 41340 48346 41368 48622
rect 41420 48612 41472 48618
rect 41420 48554 41472 48560
rect 41328 48340 41380 48346
rect 41328 48282 41380 48288
rect 41328 48068 41380 48074
rect 41328 48010 41380 48016
rect 41340 47530 41368 48010
rect 41432 47666 41460 48554
rect 41512 48204 41564 48210
rect 41512 48146 41564 48152
rect 41420 47660 41472 47666
rect 41420 47602 41472 47608
rect 41328 47524 41380 47530
rect 41328 47466 41380 47472
rect 41420 45484 41472 45490
rect 41420 45426 41472 45432
rect 41432 44878 41460 45426
rect 41524 45354 41552 48146
rect 41616 48074 41644 48690
rect 41708 48210 41736 49166
rect 41788 48680 41840 48686
rect 41788 48622 41840 48628
rect 41800 48278 41828 48622
rect 41892 48346 41920 50254
rect 41972 50176 42024 50182
rect 41972 50118 42024 50124
rect 41984 49230 42012 50118
rect 42444 49842 42472 50254
rect 43088 50182 43116 54606
rect 43180 54602 43208 55218
rect 43168 54596 43220 54602
rect 43168 54538 43220 54544
rect 43180 53650 43208 54538
rect 43548 53786 43576 56306
rect 43904 56296 43956 56302
rect 43904 56238 43956 56244
rect 43916 55418 43944 56238
rect 45192 55752 45244 55758
rect 45192 55694 45244 55700
rect 43904 55412 43956 55418
rect 43904 55354 43956 55360
rect 45008 54664 45060 54670
rect 45008 54606 45060 54612
rect 43628 54528 43680 54534
rect 43628 54470 43680 54476
rect 43640 54194 43668 54470
rect 43628 54188 43680 54194
rect 43628 54130 43680 54136
rect 43720 54188 43772 54194
rect 43720 54130 43772 54136
rect 43732 53786 43760 54130
rect 43536 53780 43588 53786
rect 43536 53722 43588 53728
rect 43720 53780 43772 53786
rect 43720 53722 43772 53728
rect 43168 53644 43220 53650
rect 43168 53586 43220 53592
rect 43720 53576 43772 53582
rect 43720 53518 43772 53524
rect 43352 53168 43404 53174
rect 43352 53110 43404 53116
rect 43364 52018 43392 53110
rect 43732 52698 43760 53518
rect 45020 53514 45048 54606
rect 45204 54330 45232 55694
rect 45388 54874 45416 56782
rect 45836 56364 45888 56370
rect 45836 56306 45888 56312
rect 45848 55962 45876 56306
rect 46572 56160 46624 56166
rect 46572 56102 46624 56108
rect 45836 55956 45888 55962
rect 45836 55898 45888 55904
rect 46584 55826 46612 56102
rect 46860 55962 46888 56782
rect 46848 55956 46900 55962
rect 46848 55898 46900 55904
rect 46940 55956 46992 55962
rect 46940 55898 46992 55904
rect 46572 55820 46624 55826
rect 46572 55762 46624 55768
rect 46952 55758 46980 55898
rect 46940 55752 46992 55758
rect 46940 55694 46992 55700
rect 45836 55276 45888 55282
rect 45836 55218 45888 55224
rect 45744 55072 45796 55078
rect 45744 55014 45796 55020
rect 45376 54868 45428 54874
rect 45376 54810 45428 54816
rect 45756 54738 45784 55014
rect 45744 54732 45796 54738
rect 45744 54674 45796 54680
rect 45652 54596 45704 54602
rect 45652 54538 45704 54544
rect 45664 54330 45692 54538
rect 45192 54324 45244 54330
rect 45192 54266 45244 54272
rect 45652 54324 45704 54330
rect 45652 54266 45704 54272
rect 45468 53984 45520 53990
rect 45468 53926 45520 53932
rect 45560 53984 45612 53990
rect 45560 53926 45612 53932
rect 45192 53644 45244 53650
rect 45192 53586 45244 53592
rect 45008 53508 45060 53514
rect 45008 53450 45060 53456
rect 44180 53100 44232 53106
rect 44180 53042 44232 53048
rect 43720 52692 43772 52698
rect 43720 52634 43772 52640
rect 43628 52420 43680 52426
rect 43628 52362 43680 52368
rect 43352 52012 43404 52018
rect 43352 51954 43404 51960
rect 43640 51406 43668 52362
rect 44192 52358 44220 53042
rect 44180 52352 44232 52358
rect 44180 52294 44232 52300
rect 43720 52012 43772 52018
rect 43772 51972 43852 52000
rect 43720 51954 43772 51960
rect 43824 51406 43852 51972
rect 43996 51944 44048 51950
rect 43996 51886 44048 51892
rect 44088 51944 44140 51950
rect 44088 51886 44140 51892
rect 43904 51468 43956 51474
rect 43904 51410 43956 51416
rect 43628 51400 43680 51406
rect 43628 51342 43680 51348
rect 43812 51400 43864 51406
rect 43812 51342 43864 51348
rect 43168 51264 43220 51270
rect 43168 51206 43220 51212
rect 43076 50176 43128 50182
rect 43076 50118 43128 50124
rect 42432 49836 42484 49842
rect 42432 49778 42484 49784
rect 42064 49632 42116 49638
rect 42064 49574 42116 49580
rect 42616 49632 42668 49638
rect 42616 49574 42668 49580
rect 41972 49224 42024 49230
rect 41972 49166 42024 49172
rect 41880 48340 41932 48346
rect 41880 48282 41932 48288
rect 41788 48272 41840 48278
rect 41788 48214 41840 48220
rect 41696 48204 41748 48210
rect 41696 48146 41748 48152
rect 41604 48068 41656 48074
rect 41604 48010 41656 48016
rect 41788 47456 41840 47462
rect 41788 47398 41840 47404
rect 41696 47184 41748 47190
rect 41696 47126 41748 47132
rect 41708 46578 41736 47126
rect 41696 46572 41748 46578
rect 41696 46514 41748 46520
rect 41512 45348 41564 45354
rect 41512 45290 41564 45296
rect 41800 44878 41828 47398
rect 42076 46646 42104 49574
rect 42628 49366 42656 49574
rect 42616 49360 42668 49366
rect 42616 49302 42668 49308
rect 42628 48890 42656 49302
rect 42616 48884 42668 48890
rect 42616 48826 42668 48832
rect 43180 48822 43208 51206
rect 43640 50930 43668 51342
rect 43916 51270 43944 51410
rect 44008 51406 44036 51886
rect 44100 51406 44128 51886
rect 43996 51400 44048 51406
rect 43996 51342 44048 51348
rect 44088 51400 44140 51406
rect 44088 51342 44140 51348
rect 43812 51264 43864 51270
rect 43812 51206 43864 51212
rect 43904 51264 43956 51270
rect 43904 51206 43956 51212
rect 43824 51074 43852 51206
rect 43824 51046 44036 51074
rect 43902 50960 43958 50969
rect 43628 50924 43680 50930
rect 43902 50895 43904 50904
rect 43628 50866 43680 50872
rect 43956 50895 43958 50904
rect 43904 50866 43956 50872
rect 44008 50862 44036 51046
rect 44100 50930 44128 51342
rect 44088 50924 44140 50930
rect 44088 50866 44140 50872
rect 43996 50856 44048 50862
rect 43996 50798 44048 50804
rect 43444 50720 43496 50726
rect 43444 50662 43496 50668
rect 43456 50454 43484 50662
rect 43444 50448 43496 50454
rect 43444 50390 43496 50396
rect 44088 50244 44140 50250
rect 44088 50186 44140 50192
rect 43444 49904 43496 49910
rect 43444 49846 43496 49852
rect 43456 49230 43484 49846
rect 43536 49632 43588 49638
rect 43536 49574 43588 49580
rect 43548 49434 43576 49574
rect 43536 49428 43588 49434
rect 43536 49370 43588 49376
rect 43444 49224 43496 49230
rect 43904 49224 43956 49230
rect 43444 49166 43496 49172
rect 43718 49192 43774 49201
rect 43904 49166 43956 49172
rect 43718 49127 43774 49136
rect 43168 48816 43220 48822
rect 43220 48764 43300 48770
rect 43168 48758 43300 48764
rect 42984 48748 43036 48754
rect 43180 48742 43300 48758
rect 43732 48754 43760 49127
rect 43916 48890 43944 49166
rect 43904 48884 43956 48890
rect 43904 48826 43956 48832
rect 42984 48690 43036 48696
rect 42996 48056 43024 48690
rect 43076 48680 43128 48686
rect 43128 48640 43208 48668
rect 43076 48622 43128 48628
rect 43180 48278 43208 48640
rect 43168 48272 43220 48278
rect 43168 48214 43220 48220
rect 43076 48068 43128 48074
rect 42996 48028 43076 48056
rect 43076 48010 43128 48016
rect 42616 48000 42668 48006
rect 42616 47942 42668 47948
rect 42628 47734 42656 47942
rect 42616 47728 42668 47734
rect 42616 47670 42668 47676
rect 42628 46714 42656 47670
rect 43088 47598 43116 48010
rect 43076 47592 43128 47598
rect 43076 47534 43128 47540
rect 43180 47462 43208 48214
rect 43272 48210 43300 48742
rect 43720 48748 43772 48754
rect 43720 48690 43772 48696
rect 43732 48346 43760 48690
rect 43720 48340 43772 48346
rect 43720 48282 43772 48288
rect 43904 48340 43956 48346
rect 43904 48282 43956 48288
rect 43260 48204 43312 48210
rect 43260 48146 43312 48152
rect 43272 47734 43300 48146
rect 43260 47728 43312 47734
rect 43260 47670 43312 47676
rect 43628 47592 43680 47598
rect 43628 47534 43680 47540
rect 43168 47456 43220 47462
rect 43168 47398 43220 47404
rect 43180 46714 43208 47398
rect 43444 46980 43496 46986
rect 43444 46922 43496 46928
rect 42616 46708 42668 46714
rect 42616 46650 42668 46656
rect 43168 46708 43220 46714
rect 43168 46650 43220 46656
rect 42064 46640 42116 46646
rect 42064 46582 42116 46588
rect 42432 46572 42484 46578
rect 42432 46514 42484 46520
rect 42156 46368 42208 46374
rect 42156 46310 42208 46316
rect 42168 45966 42196 46310
rect 42444 46170 42472 46514
rect 43456 46442 43484 46922
rect 43444 46436 43496 46442
rect 43444 46378 43496 46384
rect 43536 46436 43588 46442
rect 43536 46378 43588 46384
rect 43456 46170 43484 46378
rect 42432 46164 42484 46170
rect 42432 46106 42484 46112
rect 43444 46164 43496 46170
rect 43444 46106 43496 46112
rect 42064 45960 42116 45966
rect 42064 45902 42116 45908
rect 42156 45960 42208 45966
rect 42156 45902 42208 45908
rect 42076 45626 42104 45902
rect 42064 45620 42116 45626
rect 42064 45562 42116 45568
rect 41420 44872 41472 44878
rect 41420 44814 41472 44820
rect 41696 44872 41748 44878
rect 41696 44814 41748 44820
rect 41788 44872 41840 44878
rect 41788 44814 41840 44820
rect 41052 44464 41104 44470
rect 41052 44406 41104 44412
rect 41432 44402 41460 44814
rect 41708 44538 41736 44814
rect 43548 44810 43576 46378
rect 43640 45558 43668 47534
rect 43916 46578 43944 48282
rect 43904 46572 43956 46578
rect 43904 46514 43956 46520
rect 43628 45552 43680 45558
rect 43628 45494 43680 45500
rect 43536 44804 43588 44810
rect 43536 44746 43588 44752
rect 43812 44736 43864 44742
rect 43812 44678 43864 44684
rect 41696 44532 41748 44538
rect 41696 44474 41748 44480
rect 43824 44402 43852 44678
rect 41420 44396 41472 44402
rect 41420 44338 41472 44344
rect 42524 44396 42576 44402
rect 42524 44338 42576 44344
rect 43812 44396 43864 44402
rect 43812 44338 43864 44344
rect 42432 44260 42484 44266
rect 42432 44202 42484 44208
rect 42444 43790 42472 44202
rect 40500 43784 40552 43790
rect 40500 43726 40552 43732
rect 42432 43784 42484 43790
rect 42432 43726 42484 43732
rect 40512 43382 40540 43726
rect 42536 43722 42564 44338
rect 43168 44328 43220 44334
rect 43168 44270 43220 44276
rect 43180 43994 43208 44270
rect 43168 43988 43220 43994
rect 43168 43930 43220 43936
rect 42524 43716 42576 43722
rect 42524 43658 42576 43664
rect 40500 43376 40552 43382
rect 40500 43318 40552 43324
rect 42536 43314 42564 43658
rect 42524 43308 42576 43314
rect 42524 43250 42576 43256
rect 40960 43172 41012 43178
rect 40960 43114 41012 43120
rect 40132 42696 40184 42702
rect 40132 42638 40184 42644
rect 40316 42696 40368 42702
rect 40316 42638 40368 42644
rect 39868 41386 39988 41414
rect 39396 40520 39448 40526
rect 39396 40462 39448 40468
rect 39212 40112 39264 40118
rect 39212 40054 39264 40060
rect 39120 39840 39172 39846
rect 39040 39800 39120 39828
rect 39120 39782 39172 39788
rect 38844 39500 38896 39506
rect 38844 39442 38896 39448
rect 38752 39432 38804 39438
rect 38752 39374 38804 39380
rect 38568 38004 38620 38010
rect 38568 37946 38620 37952
rect 38752 37936 38804 37942
rect 38750 37904 38752 37913
rect 38804 37904 38806 37913
rect 39008 37868 39060 37874
rect 38750 37839 38806 37848
rect 38948 37828 39008 37856
rect 38948 37670 38976 37828
rect 39008 37810 39060 37816
rect 39028 37732 39080 37738
rect 39028 37674 39080 37680
rect 38936 37664 38988 37670
rect 38936 37606 38988 37612
rect 39040 37262 39068 37674
rect 39132 37330 39160 39782
rect 39304 37800 39356 37806
rect 39304 37742 39356 37748
rect 39316 37466 39344 37742
rect 39304 37460 39356 37466
rect 39304 37402 39356 37408
rect 39120 37324 39172 37330
rect 39120 37266 39172 37272
rect 39408 37262 39436 40462
rect 39764 40452 39816 40458
rect 39764 40394 39816 40400
rect 39580 40112 39632 40118
rect 39580 40054 39632 40060
rect 39488 39432 39540 39438
rect 39488 39374 39540 39380
rect 39500 37874 39528 39374
rect 39488 37868 39540 37874
rect 39488 37810 39540 37816
rect 39500 37466 39528 37810
rect 39488 37460 39540 37466
rect 39488 37402 39540 37408
rect 39592 37330 39620 40054
rect 39580 37324 39632 37330
rect 39580 37266 39632 37272
rect 38936 37256 38988 37262
rect 38936 37198 38988 37204
rect 39028 37256 39080 37262
rect 39028 37198 39080 37204
rect 39396 37256 39448 37262
rect 39396 37198 39448 37204
rect 39488 37256 39540 37262
rect 39488 37198 39540 37204
rect 38948 36922 38976 37198
rect 38936 36916 38988 36922
rect 38936 36858 38988 36864
rect 39028 36780 39080 36786
rect 39028 36722 39080 36728
rect 39212 36780 39264 36786
rect 39212 36722 39264 36728
rect 39040 36242 39068 36722
rect 39224 36378 39252 36722
rect 39212 36372 39264 36378
rect 39212 36314 39264 36320
rect 39028 36236 39080 36242
rect 39028 36178 39080 36184
rect 38936 36100 38988 36106
rect 38936 36042 38988 36048
rect 38948 35290 38976 36042
rect 38936 35284 38988 35290
rect 38936 35226 38988 35232
rect 39040 35170 39068 36178
rect 39224 35698 39252 36314
rect 39212 35692 39264 35698
rect 39212 35634 39264 35640
rect 39120 35488 39172 35494
rect 39120 35430 39172 35436
rect 38856 35142 39068 35170
rect 38856 33590 38884 35142
rect 39132 35086 39160 35430
rect 38936 35080 38988 35086
rect 38936 35022 38988 35028
rect 39120 35080 39172 35086
rect 39120 35022 39172 35028
rect 38948 33590 38976 35022
rect 39408 34542 39436 37198
rect 39500 34610 39528 37198
rect 39776 36174 39804 40394
rect 39868 39438 39896 41386
rect 40144 41070 40172 42638
rect 40132 41064 40184 41070
rect 40132 41006 40184 41012
rect 40314 41032 40370 41041
rect 39948 39976 40000 39982
rect 39948 39918 40000 39924
rect 39960 39642 39988 39918
rect 39948 39636 40000 39642
rect 39948 39578 40000 39584
rect 40040 39500 40092 39506
rect 40040 39442 40092 39448
rect 39856 39432 39908 39438
rect 39856 39374 39908 39380
rect 39856 39024 39908 39030
rect 39856 38966 39908 38972
rect 39868 38554 39896 38966
rect 39856 38548 39908 38554
rect 39856 38490 39908 38496
rect 39868 37874 39896 38490
rect 39948 37936 40000 37942
rect 39946 37904 39948 37913
rect 40000 37904 40002 37913
rect 39856 37868 39908 37874
rect 39946 37839 40002 37848
rect 39856 37810 39908 37816
rect 39856 37732 39908 37738
rect 40052 37720 40080 39442
rect 39908 37692 40080 37720
rect 39856 37674 39908 37680
rect 39764 36168 39816 36174
rect 39764 36110 39816 36116
rect 40052 35034 40080 37692
rect 40144 35154 40172 41006
rect 40972 41002 41000 43114
rect 41788 43104 41840 43110
rect 41788 43046 41840 43052
rect 43812 43104 43864 43110
rect 43812 43046 43864 43052
rect 41800 42702 41828 43046
rect 41788 42696 41840 42702
rect 41788 42638 41840 42644
rect 41880 42696 41932 42702
rect 41880 42638 41932 42644
rect 43352 42696 43404 42702
rect 43352 42638 43404 42644
rect 41328 42560 41380 42566
rect 41328 42502 41380 42508
rect 41340 42226 41368 42502
rect 41892 42294 41920 42638
rect 43364 42294 43392 42638
rect 41880 42288 41932 42294
rect 41880 42230 41932 42236
rect 43352 42288 43404 42294
rect 43352 42230 43404 42236
rect 43824 42226 43852 43046
rect 44100 42634 44128 50186
rect 44192 49706 44220 52294
rect 45204 51406 45232 53586
rect 45480 52426 45508 53926
rect 45572 53242 45600 53926
rect 45848 53786 45876 55218
rect 46952 54874 46980 55694
rect 46940 54868 46992 54874
rect 46940 54810 46992 54816
rect 46572 54528 46624 54534
rect 46572 54470 46624 54476
rect 46584 54126 46612 54470
rect 46952 54194 46980 54810
rect 46940 54188 46992 54194
rect 46940 54130 46992 54136
rect 46572 54120 46624 54126
rect 46572 54062 46624 54068
rect 45836 53780 45888 53786
rect 45836 53722 45888 53728
rect 46584 53650 46612 54062
rect 46572 53644 46624 53650
rect 46572 53586 46624 53592
rect 46112 53576 46164 53582
rect 46112 53518 46164 53524
rect 45560 53236 45612 53242
rect 45560 53178 45612 53184
rect 45652 53100 45704 53106
rect 45652 53042 45704 53048
rect 45560 52556 45612 52562
rect 45560 52498 45612 52504
rect 45572 52426 45600 52498
rect 45468 52420 45520 52426
rect 45468 52362 45520 52368
rect 45560 52420 45612 52426
rect 45560 52362 45612 52368
rect 45664 52018 45692 53042
rect 46124 53038 46152 53518
rect 46204 53440 46256 53446
rect 46204 53382 46256 53388
rect 46388 53440 46440 53446
rect 46388 53382 46440 53388
rect 46216 53106 46244 53382
rect 46400 53174 46428 53382
rect 46388 53168 46440 53174
rect 46388 53110 46440 53116
rect 46204 53100 46256 53106
rect 46204 53042 46256 53048
rect 46112 53032 46164 53038
rect 46112 52974 46164 52980
rect 45744 52624 45796 52630
rect 45744 52566 45796 52572
rect 45652 52012 45704 52018
rect 45652 51954 45704 51960
rect 45192 51400 45244 51406
rect 45192 51342 45244 51348
rect 45468 51400 45520 51406
rect 45468 51342 45520 51348
rect 44640 49904 44692 49910
rect 44640 49846 44692 49852
rect 44180 49700 44232 49706
rect 44180 49642 44232 49648
rect 44272 48136 44324 48142
rect 44272 48078 44324 48084
rect 44456 48136 44508 48142
rect 44456 48078 44508 48084
rect 44284 47598 44312 48078
rect 44272 47592 44324 47598
rect 44272 47534 44324 47540
rect 44364 47456 44416 47462
rect 44364 47398 44416 47404
rect 44376 47258 44404 47398
rect 44364 47252 44416 47258
rect 44364 47194 44416 47200
rect 44376 46578 44404 47194
rect 44468 47054 44496 48078
rect 44652 47530 44680 49846
rect 44916 49836 44968 49842
rect 44916 49778 44968 49784
rect 45008 49836 45060 49842
rect 45008 49778 45060 49784
rect 44928 49638 44956 49778
rect 44916 49632 44968 49638
rect 44916 49574 44968 49580
rect 45020 48210 45048 49778
rect 45100 49700 45152 49706
rect 45100 49642 45152 49648
rect 45112 49162 45140 49642
rect 45376 49632 45428 49638
rect 45376 49574 45428 49580
rect 45388 49230 45416 49574
rect 45376 49224 45428 49230
rect 45376 49166 45428 49172
rect 45100 49156 45152 49162
rect 45100 49098 45152 49104
rect 45112 48754 45140 49098
rect 45376 49088 45428 49094
rect 45376 49030 45428 49036
rect 45100 48748 45152 48754
rect 45100 48690 45152 48696
rect 45192 48544 45244 48550
rect 45192 48486 45244 48492
rect 45008 48204 45060 48210
rect 45008 48146 45060 48152
rect 44916 48136 44968 48142
rect 44916 48078 44968 48084
rect 44928 47666 44956 48078
rect 44916 47660 44968 47666
rect 44916 47602 44968 47608
rect 44640 47524 44692 47530
rect 44640 47466 44692 47472
rect 44928 47054 44956 47602
rect 45204 47462 45232 48486
rect 45388 48314 45416 49030
rect 45296 48286 45416 48314
rect 45296 48142 45324 48286
rect 45480 48142 45508 51342
rect 45664 51338 45692 51954
rect 45652 51332 45704 51338
rect 45652 51274 45704 51280
rect 45664 50930 45692 51274
rect 45652 50924 45704 50930
rect 45652 50866 45704 50872
rect 45664 50250 45692 50866
rect 45652 50244 45704 50250
rect 45652 50186 45704 50192
rect 45652 49768 45704 49774
rect 45652 49710 45704 49716
rect 45560 49360 45612 49366
rect 45560 49302 45612 49308
rect 45284 48136 45336 48142
rect 45284 48078 45336 48084
rect 45468 48136 45520 48142
rect 45468 48078 45520 48084
rect 45192 47456 45244 47462
rect 45192 47398 45244 47404
rect 44456 47048 44508 47054
rect 44456 46990 44508 46996
rect 44916 47048 44968 47054
rect 44916 46990 44968 46996
rect 44364 46572 44416 46578
rect 44364 46514 44416 46520
rect 45100 46368 45152 46374
rect 45100 46310 45152 46316
rect 45112 46102 45140 46310
rect 45296 46170 45324 48078
rect 45572 46714 45600 49302
rect 45664 49230 45692 49710
rect 45652 49224 45704 49230
rect 45650 49192 45652 49201
rect 45704 49192 45706 49201
rect 45650 49127 45706 49136
rect 45756 48822 45784 52566
rect 46124 52494 46152 52974
rect 46216 52698 46244 53042
rect 46296 52896 46348 52902
rect 46296 52838 46348 52844
rect 46204 52692 46256 52698
rect 46204 52634 46256 52640
rect 46112 52488 46164 52494
rect 46112 52430 46164 52436
rect 46124 51406 46152 52430
rect 46308 52018 46336 52838
rect 46296 52012 46348 52018
rect 46296 51954 46348 51960
rect 46400 51898 46428 53110
rect 46584 52494 46612 53586
rect 46940 53168 46992 53174
rect 46940 53110 46992 53116
rect 46572 52488 46624 52494
rect 46572 52430 46624 52436
rect 46480 52012 46532 52018
rect 46480 51954 46532 51960
rect 46308 51882 46428 51898
rect 46296 51876 46428 51882
rect 46348 51870 46428 51876
rect 46296 51818 46348 51824
rect 46112 51400 46164 51406
rect 46112 51342 46164 51348
rect 45836 51264 45888 51270
rect 45836 51206 45888 51212
rect 45848 50318 45876 51206
rect 46308 50998 46336 51818
rect 46492 51074 46520 51954
rect 46584 51406 46612 52430
rect 46952 52358 46980 53110
rect 46940 52352 46992 52358
rect 46940 52294 46992 52300
rect 46572 51400 46624 51406
rect 46572 51342 46624 51348
rect 46388 51060 46440 51066
rect 46492 51046 46612 51074
rect 46388 51002 46440 51008
rect 46296 50992 46348 50998
rect 46296 50934 46348 50940
rect 46204 50788 46256 50794
rect 46204 50730 46256 50736
rect 45836 50312 45888 50318
rect 45836 50254 45888 50260
rect 45928 50176 45980 50182
rect 45928 50118 45980 50124
rect 46112 50176 46164 50182
rect 46112 50118 46164 50124
rect 45940 49978 45968 50118
rect 45928 49972 45980 49978
rect 45928 49914 45980 49920
rect 45928 49088 45980 49094
rect 45928 49030 45980 49036
rect 45940 48890 45968 49030
rect 45928 48884 45980 48890
rect 45928 48826 45980 48832
rect 46020 48884 46072 48890
rect 46020 48826 46072 48832
rect 45744 48816 45796 48822
rect 45744 48758 45796 48764
rect 45652 48612 45704 48618
rect 45652 48554 45704 48560
rect 45664 48074 45692 48554
rect 46032 48346 46060 48826
rect 46020 48340 46072 48346
rect 46020 48282 46072 48288
rect 45652 48068 45704 48074
rect 45652 48010 45704 48016
rect 45652 47660 45704 47666
rect 45652 47602 45704 47608
rect 45664 47054 45692 47602
rect 46124 47258 46152 50118
rect 46216 48754 46244 50730
rect 46296 50312 46348 50318
rect 46296 50254 46348 50260
rect 46308 49774 46336 50254
rect 46400 49978 46428 51002
rect 46388 49972 46440 49978
rect 46388 49914 46440 49920
rect 46296 49768 46348 49774
rect 46296 49710 46348 49716
rect 46308 49434 46336 49710
rect 46480 49632 46532 49638
rect 46480 49574 46532 49580
rect 46296 49428 46348 49434
rect 46296 49370 46348 49376
rect 46492 49230 46520 49574
rect 46480 49224 46532 49230
rect 46480 49166 46532 49172
rect 46204 48748 46256 48754
rect 46204 48690 46256 48696
rect 46216 48550 46244 48690
rect 46204 48544 46256 48550
rect 46204 48486 46256 48492
rect 46296 47592 46348 47598
rect 46296 47534 46348 47540
rect 46308 47258 46336 47534
rect 46112 47252 46164 47258
rect 46112 47194 46164 47200
rect 46296 47252 46348 47258
rect 46296 47194 46348 47200
rect 45836 47116 45888 47122
rect 45836 47058 45888 47064
rect 45652 47048 45704 47054
rect 45652 46990 45704 46996
rect 45560 46708 45612 46714
rect 45560 46650 45612 46656
rect 45664 46578 45692 46990
rect 45652 46572 45704 46578
rect 45652 46514 45704 46520
rect 45664 46170 45692 46514
rect 45848 46510 45876 47058
rect 45836 46504 45888 46510
rect 45836 46446 45888 46452
rect 45284 46164 45336 46170
rect 45284 46106 45336 46112
rect 45652 46164 45704 46170
rect 45652 46106 45704 46112
rect 45100 46096 45152 46102
rect 45100 46038 45152 46044
rect 45848 45898 45876 46446
rect 45836 45892 45888 45898
rect 45836 45834 45888 45840
rect 44916 45484 44968 45490
rect 44916 45426 44968 45432
rect 45652 45484 45704 45490
rect 45652 45426 45704 45432
rect 44180 44940 44232 44946
rect 44180 44882 44232 44888
rect 44192 44742 44220 44882
rect 44364 44872 44416 44878
rect 44364 44814 44416 44820
rect 44180 44736 44232 44742
rect 44180 44678 44232 44684
rect 44192 43790 44220 44678
rect 44376 43994 44404 44814
rect 44928 44538 44956 45426
rect 45560 45280 45612 45286
rect 45560 45222 45612 45228
rect 45572 45082 45600 45222
rect 45560 45076 45612 45082
rect 45560 45018 45612 45024
rect 44916 44532 44968 44538
rect 44916 44474 44968 44480
rect 44364 43988 44416 43994
rect 44364 43930 44416 43936
rect 44928 43858 44956 44474
rect 45572 44198 45600 45018
rect 45664 44878 45692 45426
rect 45744 45416 45796 45422
rect 45744 45358 45796 45364
rect 45756 44946 45784 45358
rect 45744 44940 45796 44946
rect 45744 44882 45796 44888
rect 45652 44872 45704 44878
rect 45652 44814 45704 44820
rect 45756 44402 45784 44882
rect 45848 44538 45876 45834
rect 46308 45014 46336 47194
rect 46388 47048 46440 47054
rect 46388 46990 46440 46996
rect 46400 46918 46428 46990
rect 46388 46912 46440 46918
rect 46388 46854 46440 46860
rect 46400 45966 46428 46854
rect 46388 45960 46440 45966
rect 46388 45902 46440 45908
rect 46296 45008 46348 45014
rect 46296 44950 46348 44956
rect 46204 44872 46256 44878
rect 46204 44814 46256 44820
rect 45836 44532 45888 44538
rect 45836 44474 45888 44480
rect 45744 44396 45796 44402
rect 45744 44338 45796 44344
rect 45652 44260 45704 44266
rect 45652 44202 45704 44208
rect 45560 44192 45612 44198
rect 45560 44134 45612 44140
rect 45664 43858 45692 44202
rect 44916 43852 44968 43858
rect 44916 43794 44968 43800
rect 45652 43852 45704 43858
rect 45652 43794 45704 43800
rect 44180 43784 44232 43790
rect 45756 43738 45784 44338
rect 46216 44334 46244 44814
rect 46204 44328 46256 44334
rect 46204 44270 46256 44276
rect 46216 43790 46244 44270
rect 44180 43726 44232 43732
rect 44192 43246 44220 43726
rect 45664 43710 45784 43738
rect 46204 43784 46256 43790
rect 46204 43726 46256 43732
rect 46388 43716 46440 43722
rect 45664 43654 45692 43710
rect 46388 43658 46440 43664
rect 45652 43648 45704 43654
rect 45652 43590 45704 43596
rect 45664 43314 45692 43590
rect 46400 43450 46428 43658
rect 46388 43444 46440 43450
rect 46388 43386 46440 43392
rect 45652 43308 45704 43314
rect 45652 43250 45704 43256
rect 44180 43240 44232 43246
rect 44180 43182 44232 43188
rect 46584 42770 46612 51046
rect 46664 51060 46716 51066
rect 46664 51002 46716 51008
rect 46676 47258 46704 51002
rect 46952 48890 46980 52294
rect 47032 50856 47084 50862
rect 47032 50798 47084 50804
rect 47044 50522 47072 50798
rect 47124 50788 47176 50794
rect 47124 50730 47176 50736
rect 47032 50516 47084 50522
rect 47032 50458 47084 50464
rect 47136 50386 47164 50730
rect 47308 50720 47360 50726
rect 47308 50662 47360 50668
rect 47320 50522 47348 50662
rect 47308 50516 47360 50522
rect 47308 50458 47360 50464
rect 47124 50380 47176 50386
rect 47124 50322 47176 50328
rect 46940 48884 46992 48890
rect 46940 48826 46992 48832
rect 47032 48544 47084 48550
rect 47032 48486 47084 48492
rect 47044 48278 47072 48486
rect 47032 48272 47084 48278
rect 47032 48214 47084 48220
rect 47124 48204 47176 48210
rect 47124 48146 47176 48152
rect 46664 47252 46716 47258
rect 46664 47194 46716 47200
rect 47136 46646 47164 48146
rect 47216 48000 47268 48006
rect 47216 47942 47268 47948
rect 47228 46646 47256 47942
rect 47124 46640 47176 46646
rect 47124 46582 47176 46588
rect 47216 46640 47268 46646
rect 47216 46582 47268 46588
rect 46664 45076 46716 45082
rect 46664 45018 46716 45024
rect 46676 44742 46704 45018
rect 46664 44736 46716 44742
rect 46664 44678 46716 44684
rect 46572 42764 46624 42770
rect 46572 42706 46624 42712
rect 44088 42628 44140 42634
rect 44088 42570 44140 42576
rect 45284 42628 45336 42634
rect 45284 42570 45336 42576
rect 45008 42560 45060 42566
rect 45008 42502 45060 42508
rect 45020 42294 45048 42502
rect 45008 42288 45060 42294
rect 45008 42230 45060 42236
rect 41328 42220 41380 42226
rect 41328 42162 41380 42168
rect 41696 42220 41748 42226
rect 41696 42162 41748 42168
rect 43628 42220 43680 42226
rect 43812 42220 43864 42226
rect 43680 42180 43760 42208
rect 43628 42162 43680 42168
rect 41340 41614 41368 42162
rect 41328 41608 41380 41614
rect 41328 41550 41380 41556
rect 41432 41546 41552 41562
rect 41432 41540 41564 41546
rect 41432 41534 41512 41540
rect 40314 40967 40370 40976
rect 40960 40996 41012 41002
rect 40328 40934 40356 40967
rect 40960 40938 41012 40944
rect 40316 40928 40368 40934
rect 40316 40870 40368 40876
rect 40500 40044 40552 40050
rect 40500 39986 40552 39992
rect 40512 39098 40540 39986
rect 40868 39432 40920 39438
rect 40972 39420 41000 40938
rect 41432 40662 41460 41534
rect 41512 41482 41564 41488
rect 41708 41414 41736 42162
rect 42432 42152 42484 42158
rect 42432 42094 42484 42100
rect 42246 41848 42302 41857
rect 42246 41783 42302 41792
rect 42260 41682 42288 41783
rect 42444 41682 42472 42094
rect 43168 42084 43220 42090
rect 43168 42026 43220 42032
rect 42248 41676 42300 41682
rect 42248 41618 42300 41624
rect 42432 41676 42484 41682
rect 42432 41618 42484 41624
rect 43180 41614 43208 42026
rect 42340 41608 42392 41614
rect 42340 41550 42392 41556
rect 43168 41608 43220 41614
rect 43168 41550 43220 41556
rect 42352 41478 42380 41550
rect 42892 41540 42944 41546
rect 42892 41482 42944 41488
rect 41972 41472 42024 41478
rect 41972 41414 42024 41420
rect 42340 41472 42392 41478
rect 42340 41414 42392 41420
rect 42800 41472 42852 41478
rect 42800 41414 42852 41420
rect 41524 41386 41736 41414
rect 41524 41070 41552 41386
rect 41512 41064 41564 41070
rect 41512 41006 41564 41012
rect 41984 40934 42012 41414
rect 42340 41268 42392 41274
rect 42340 41210 42392 41216
rect 41972 40928 42024 40934
rect 41972 40870 42024 40876
rect 41420 40656 41472 40662
rect 41420 40598 41472 40604
rect 41432 40118 41460 40598
rect 42352 40594 42380 41210
rect 42524 41200 42576 41206
rect 42524 41142 42576 41148
rect 42340 40588 42392 40594
rect 42340 40530 42392 40536
rect 42536 40458 42564 41142
rect 42812 41070 42840 41414
rect 42904 41206 42932 41482
rect 42892 41200 42944 41206
rect 42892 41142 42944 41148
rect 42616 41064 42668 41070
rect 42616 41006 42668 41012
rect 42800 41064 42852 41070
rect 42800 41006 42852 41012
rect 42892 41064 42944 41070
rect 42892 41006 42944 41012
rect 42628 40730 42656 41006
rect 42616 40724 42668 40730
rect 42616 40666 42668 40672
rect 42524 40452 42576 40458
rect 42524 40394 42576 40400
rect 42536 40118 42564 40394
rect 41420 40112 41472 40118
rect 41420 40054 41472 40060
rect 42524 40112 42576 40118
rect 42524 40054 42576 40060
rect 41052 39840 41104 39846
rect 41052 39782 41104 39788
rect 41064 39438 41092 39782
rect 40920 39392 41000 39420
rect 40868 39374 40920 39380
rect 40684 39296 40736 39302
rect 40684 39238 40736 39244
rect 40500 39092 40552 39098
rect 40500 39034 40552 39040
rect 40696 38962 40724 39238
rect 40684 38956 40736 38962
rect 40684 38898 40736 38904
rect 40972 38350 41000 39392
rect 41052 39432 41104 39438
rect 41052 39374 41104 39380
rect 41064 39030 41092 39374
rect 41052 39024 41104 39030
rect 41052 38966 41104 38972
rect 41432 38962 41460 40054
rect 42616 39840 42668 39846
rect 42616 39782 42668 39788
rect 42628 39438 42656 39782
rect 42812 39438 42840 41006
rect 42904 39506 42932 41006
rect 43628 40928 43680 40934
rect 43628 40870 43680 40876
rect 43352 40112 43404 40118
rect 43352 40054 43404 40060
rect 42892 39500 42944 39506
rect 42892 39442 42944 39448
rect 42616 39432 42668 39438
rect 42616 39374 42668 39380
rect 42800 39432 42852 39438
rect 42800 39374 42852 39380
rect 42340 39364 42392 39370
rect 42340 39306 42392 39312
rect 42524 39364 42576 39370
rect 42524 39306 42576 39312
rect 42352 38962 42380 39306
rect 42536 39098 42564 39306
rect 42524 39092 42576 39098
rect 42524 39034 42576 39040
rect 41420 38956 41472 38962
rect 41420 38898 41472 38904
rect 42340 38956 42392 38962
rect 42340 38898 42392 38904
rect 42812 38894 42840 39374
rect 42904 38962 42932 39442
rect 43260 39296 43312 39302
rect 43260 39238 43312 39244
rect 43272 39030 43300 39238
rect 43260 39024 43312 39030
rect 43260 38966 43312 38972
rect 43364 38962 43392 40054
rect 43640 40050 43668 40870
rect 43732 40526 43760 42180
rect 43812 42162 43864 42168
rect 43904 41132 43956 41138
rect 43904 41074 43956 41080
rect 43916 40730 43944 41074
rect 44180 40928 44232 40934
rect 44180 40870 44232 40876
rect 43904 40724 43956 40730
rect 43904 40666 43956 40672
rect 43720 40520 43772 40526
rect 43720 40462 43772 40468
rect 43628 40044 43680 40050
rect 43628 39986 43680 39992
rect 43444 39296 43496 39302
rect 43444 39238 43496 39244
rect 42892 38956 42944 38962
rect 42892 38898 42944 38904
rect 43352 38956 43404 38962
rect 43352 38898 43404 38904
rect 42800 38888 42852 38894
rect 42800 38830 42852 38836
rect 42708 38820 42760 38826
rect 42708 38762 42760 38768
rect 40960 38344 41012 38350
rect 40960 38286 41012 38292
rect 40592 38276 40644 38282
rect 40592 38218 40644 38224
rect 40604 36854 40632 38218
rect 40868 38004 40920 38010
rect 40868 37946 40920 37952
rect 40684 37460 40736 37466
rect 40684 37402 40736 37408
rect 40592 36848 40644 36854
rect 40592 36790 40644 36796
rect 40408 36576 40460 36582
rect 40408 36518 40460 36524
rect 40316 35692 40368 35698
rect 40316 35634 40368 35640
rect 40328 35154 40356 35634
rect 40132 35148 40184 35154
rect 40132 35090 40184 35096
rect 40316 35148 40368 35154
rect 40316 35090 40368 35096
rect 40052 35006 40172 35034
rect 39488 34604 39540 34610
rect 39488 34546 39540 34552
rect 39120 34536 39172 34542
rect 39120 34478 39172 34484
rect 39396 34536 39448 34542
rect 39396 34478 39448 34484
rect 39028 33856 39080 33862
rect 39028 33798 39080 33804
rect 38844 33584 38896 33590
rect 38844 33526 38896 33532
rect 38936 33584 38988 33590
rect 38936 33526 38988 33532
rect 38856 31822 38884 33526
rect 39040 33522 39068 33798
rect 39132 33658 39160 34478
rect 39120 33652 39172 33658
rect 39120 33594 39172 33600
rect 39028 33516 39080 33522
rect 39028 33458 39080 33464
rect 39304 32768 39356 32774
rect 39304 32710 39356 32716
rect 39316 32434 39344 32710
rect 39408 32502 39436 34478
rect 39500 32502 39528 34546
rect 40040 33924 40092 33930
rect 40040 33866 40092 33872
rect 40052 33658 40080 33866
rect 40040 33652 40092 33658
rect 40040 33594 40092 33600
rect 40040 33516 40092 33522
rect 40040 33458 40092 33464
rect 39396 32496 39448 32502
rect 39396 32438 39448 32444
rect 39488 32496 39540 32502
rect 39488 32438 39540 32444
rect 39304 32428 39356 32434
rect 39304 32370 39356 32376
rect 38844 31816 38896 31822
rect 38844 31758 38896 31764
rect 38856 31414 38884 31758
rect 38844 31408 38896 31414
rect 38844 31350 38896 31356
rect 39212 31408 39264 31414
rect 39212 31350 39264 31356
rect 38936 31340 38988 31346
rect 38936 31282 38988 31288
rect 38844 30592 38896 30598
rect 38948 30580 38976 31282
rect 39120 31136 39172 31142
rect 39120 31078 39172 31084
rect 38896 30552 38976 30580
rect 38844 30534 38896 30540
rect 38856 29646 38884 30534
rect 39132 30258 39160 31078
rect 39120 30252 39172 30258
rect 39120 30194 39172 30200
rect 38936 30048 38988 30054
rect 38936 29990 38988 29996
rect 38844 29640 38896 29646
rect 38844 29582 38896 29588
rect 38948 29510 38976 29990
rect 39224 29646 39252 31350
rect 39500 30258 39528 32438
rect 39580 32428 39632 32434
rect 39580 32370 39632 32376
rect 39592 31482 39620 32370
rect 40052 31822 40080 33458
rect 40144 33402 40172 35006
rect 40224 34740 40276 34746
rect 40224 34682 40276 34688
rect 40236 33590 40264 34682
rect 40328 33658 40356 35090
rect 40420 34066 40448 36518
rect 40500 35624 40552 35630
rect 40500 35566 40552 35572
rect 40512 34746 40540 35566
rect 40500 34740 40552 34746
rect 40500 34682 40552 34688
rect 40408 34060 40460 34066
rect 40408 34002 40460 34008
rect 40316 33652 40368 33658
rect 40316 33594 40368 33600
rect 40224 33584 40276 33590
rect 40224 33526 40276 33532
rect 40144 33386 40356 33402
rect 40144 33380 40368 33386
rect 40144 33374 40316 33380
rect 40316 33322 40368 33328
rect 40040 31816 40092 31822
rect 40092 31764 40172 31770
rect 40040 31758 40172 31764
rect 40052 31742 40172 31758
rect 39580 31476 39632 31482
rect 39580 31418 39632 31424
rect 40040 30728 40092 30734
rect 40040 30670 40092 30676
rect 40052 30394 40080 30670
rect 40144 30666 40172 31742
rect 40224 31680 40276 31686
rect 40224 31622 40276 31628
rect 40236 31346 40264 31622
rect 40224 31340 40276 31346
rect 40224 31282 40276 31288
rect 40132 30660 40184 30666
rect 40132 30602 40184 30608
rect 40040 30388 40092 30394
rect 40040 30330 40092 30336
rect 39488 30252 39540 30258
rect 39488 30194 39540 30200
rect 40052 29646 40080 30330
rect 39212 29640 39264 29646
rect 39212 29582 39264 29588
rect 40040 29640 40092 29646
rect 40040 29582 40092 29588
rect 40144 29578 40172 30602
rect 40328 30274 40356 33322
rect 40236 30246 40356 30274
rect 40132 29572 40184 29578
rect 40132 29514 40184 29520
rect 38936 29504 38988 29510
rect 38936 29446 38988 29452
rect 39488 29504 39540 29510
rect 39488 29446 39540 29452
rect 39500 29170 39528 29446
rect 40236 29170 40264 30246
rect 40316 30184 40368 30190
rect 40316 30126 40368 30132
rect 40328 29578 40356 30126
rect 40316 29572 40368 29578
rect 40316 29514 40368 29520
rect 39304 29164 39356 29170
rect 39304 29106 39356 29112
rect 39488 29164 39540 29170
rect 39488 29106 39540 29112
rect 40224 29164 40276 29170
rect 40224 29106 40276 29112
rect 39316 29034 39344 29106
rect 39304 29028 39356 29034
rect 39304 28970 39356 28976
rect 40224 29028 40276 29034
rect 40224 28970 40276 28976
rect 39120 28960 39172 28966
rect 39120 28902 39172 28908
rect 39132 28082 39160 28902
rect 39120 28076 39172 28082
rect 39120 28018 39172 28024
rect 40040 28076 40092 28082
rect 40040 28018 40092 28024
rect 38476 27600 38528 27606
rect 38476 27542 38528 27548
rect 37372 27396 37424 27402
rect 37372 27338 37424 27344
rect 37384 27130 37412 27338
rect 37372 27124 37424 27130
rect 37372 27066 37424 27072
rect 40052 26994 40080 28018
rect 40236 27878 40264 28970
rect 40420 28626 40448 34002
rect 40696 33522 40724 37402
rect 40880 37262 40908 37946
rect 40868 37256 40920 37262
rect 40868 37198 40920 37204
rect 40972 35018 41000 38286
rect 42720 37874 42748 38762
rect 42708 37868 42760 37874
rect 42708 37810 42760 37816
rect 41880 37256 41932 37262
rect 41880 37198 41932 37204
rect 41892 36786 41920 37198
rect 42720 36922 42748 37810
rect 42812 37262 42840 38830
rect 43456 38350 43484 39238
rect 43732 39030 43760 40462
rect 44192 40118 44220 40870
rect 45008 40588 45060 40594
rect 45008 40530 45060 40536
rect 44364 40180 44416 40186
rect 44364 40122 44416 40128
rect 44180 40112 44232 40118
rect 44180 40054 44232 40060
rect 43812 39432 43864 39438
rect 43812 39374 43864 39380
rect 43824 39098 43852 39374
rect 43812 39092 43864 39098
rect 43812 39034 43864 39040
rect 43720 39024 43772 39030
rect 43720 38966 43772 38972
rect 44088 38888 44140 38894
rect 44088 38830 44140 38836
rect 44100 38486 44128 38830
rect 44088 38480 44140 38486
rect 44088 38422 44140 38428
rect 43444 38344 43496 38350
rect 43444 38286 43496 38292
rect 44376 37942 44404 40122
rect 44916 39296 44968 39302
rect 44916 39238 44968 39244
rect 44928 38962 44956 39238
rect 44916 38956 44968 38962
rect 44916 38898 44968 38904
rect 44364 37936 44416 37942
rect 44364 37878 44416 37884
rect 43076 37392 43128 37398
rect 43076 37334 43128 37340
rect 42800 37256 42852 37262
rect 42800 37198 42852 37204
rect 42708 36916 42760 36922
rect 42708 36858 42760 36864
rect 42432 36848 42484 36854
rect 42432 36790 42484 36796
rect 41880 36780 41932 36786
rect 41880 36722 41932 36728
rect 41328 36576 41380 36582
rect 41328 36518 41380 36524
rect 41340 36378 41368 36518
rect 41328 36372 41380 36378
rect 41328 36314 41380 36320
rect 42444 36174 42472 36790
rect 42720 36718 42748 36858
rect 42708 36712 42760 36718
rect 42708 36654 42760 36660
rect 42800 36644 42852 36650
rect 42800 36586 42852 36592
rect 42432 36168 42484 36174
rect 42432 36110 42484 36116
rect 42444 35766 42472 36110
rect 42812 35766 42840 36586
rect 42984 36168 43036 36174
rect 42984 36110 43036 36116
rect 42432 35760 42484 35766
rect 42432 35702 42484 35708
rect 42800 35760 42852 35766
rect 42800 35702 42852 35708
rect 41604 35692 41656 35698
rect 41604 35634 41656 35640
rect 40960 35012 41012 35018
rect 40960 34954 41012 34960
rect 40972 34610 41000 34954
rect 41616 34746 41644 35634
rect 41788 34944 41840 34950
rect 41788 34886 41840 34892
rect 41604 34740 41656 34746
rect 41604 34682 41656 34688
rect 41800 34610 41828 34886
rect 40960 34604 41012 34610
rect 40960 34546 41012 34552
rect 41788 34604 41840 34610
rect 41788 34546 41840 34552
rect 42064 33992 42116 33998
rect 42064 33934 42116 33940
rect 41328 33924 41380 33930
rect 41328 33866 41380 33872
rect 41236 33856 41288 33862
rect 41236 33798 41288 33804
rect 40684 33516 40736 33522
rect 40684 33458 40736 33464
rect 41248 33318 41276 33798
rect 41236 33312 41288 33318
rect 41236 33254 41288 33260
rect 41144 32428 41196 32434
rect 41144 32370 41196 32376
rect 40684 32224 40736 32230
rect 40684 32166 40736 32172
rect 40696 31890 40724 32166
rect 40684 31884 40736 31890
rect 40684 31826 40736 31832
rect 41156 31754 41184 32370
rect 41144 31748 41196 31754
rect 41144 31690 41196 31696
rect 41156 30734 41184 31690
rect 41144 30728 41196 30734
rect 41144 30670 41196 30676
rect 40776 30592 40828 30598
rect 40776 30534 40828 30540
rect 40592 30252 40644 30258
rect 40592 30194 40644 30200
rect 40604 29306 40632 30194
rect 40684 29504 40736 29510
rect 40684 29446 40736 29452
rect 40592 29300 40644 29306
rect 40592 29242 40644 29248
rect 40408 28620 40460 28626
rect 40408 28562 40460 28568
rect 40420 28150 40448 28562
rect 40408 28144 40460 28150
rect 40408 28086 40460 28092
rect 40696 28014 40724 29446
rect 40788 29170 40816 30534
rect 40776 29164 40828 29170
rect 40776 29106 40828 29112
rect 40868 28484 40920 28490
rect 40868 28426 40920 28432
rect 40880 28218 40908 28426
rect 41052 28416 41104 28422
rect 41052 28358 41104 28364
rect 40868 28212 40920 28218
rect 40868 28154 40920 28160
rect 41064 28082 41092 28358
rect 41052 28076 41104 28082
rect 41052 28018 41104 28024
rect 40684 28008 40736 28014
rect 40684 27950 40736 27956
rect 40224 27872 40276 27878
rect 40224 27814 40276 27820
rect 40236 27606 40264 27814
rect 40224 27600 40276 27606
rect 40224 27542 40276 27548
rect 40868 27464 40920 27470
rect 40868 27406 40920 27412
rect 40040 26988 40092 26994
rect 40040 26930 40092 26936
rect 40316 26920 40368 26926
rect 40316 26862 40368 26868
rect 38844 26852 38896 26858
rect 38844 26794 38896 26800
rect 36912 18080 36964 18086
rect 36912 18022 36964 18028
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 38856 16574 38884 26794
rect 40328 26586 40356 26862
rect 40316 26580 40368 26586
rect 40316 26522 40368 26528
rect 40880 26450 40908 27406
rect 41248 26450 41276 33254
rect 41340 32366 41368 33866
rect 41328 32360 41380 32366
rect 41328 32302 41380 32308
rect 42076 32298 42104 33934
rect 42444 32910 42472 35702
rect 42800 35624 42852 35630
rect 42800 35566 42852 35572
rect 42812 35154 42840 35566
rect 42800 35148 42852 35154
rect 42800 35090 42852 35096
rect 42996 35086 43024 36110
rect 42984 35080 43036 35086
rect 42984 35022 43036 35028
rect 42800 34128 42852 34134
rect 42800 34070 42852 34076
rect 42812 33674 42840 34070
rect 42812 33646 42932 33674
rect 42800 33516 42852 33522
rect 42800 33458 42852 33464
rect 42812 32910 42840 33458
rect 42904 33114 42932 33646
rect 42996 33522 43024 35022
rect 43088 33998 43116 37334
rect 44376 37262 44404 37878
rect 45020 37874 45048 40530
rect 45192 40452 45244 40458
rect 45192 40394 45244 40400
rect 45204 40186 45232 40394
rect 45192 40180 45244 40186
rect 45192 40122 45244 40128
rect 45100 39432 45152 39438
rect 45100 39374 45152 39380
rect 45112 39098 45140 39374
rect 45100 39092 45152 39098
rect 45100 39034 45152 39040
rect 45192 39024 45244 39030
rect 45192 38966 45244 38972
rect 45204 38554 45232 38966
rect 45192 38548 45244 38554
rect 45192 38490 45244 38496
rect 45008 37868 45060 37874
rect 45008 37810 45060 37816
rect 44916 37664 44968 37670
rect 44916 37606 44968 37612
rect 44364 37256 44416 37262
rect 44364 37198 44416 37204
rect 43260 37188 43312 37194
rect 43260 37130 43312 37136
rect 44732 37188 44784 37194
rect 44732 37130 44784 37136
rect 44824 37188 44876 37194
rect 44824 37130 44876 37136
rect 43272 36786 43300 37130
rect 43352 36916 43404 36922
rect 43352 36858 43404 36864
rect 43260 36780 43312 36786
rect 43260 36722 43312 36728
rect 43272 34066 43300 36722
rect 43364 36718 43392 36858
rect 43352 36712 43404 36718
rect 43352 36654 43404 36660
rect 44744 36650 44772 37130
rect 44836 36922 44864 37130
rect 44928 36922 44956 37606
rect 45204 37262 45232 38490
rect 45192 37256 45244 37262
rect 45192 37198 45244 37204
rect 45008 37120 45060 37126
rect 45008 37062 45060 37068
rect 44824 36916 44876 36922
rect 44824 36858 44876 36864
rect 44916 36916 44968 36922
rect 44916 36858 44968 36864
rect 44824 36780 44876 36786
rect 44824 36722 44876 36728
rect 44732 36644 44784 36650
rect 44732 36586 44784 36592
rect 44836 36242 44864 36722
rect 44916 36712 44968 36718
rect 45020 36700 45048 37062
rect 44968 36672 45048 36700
rect 44916 36654 44968 36660
rect 45192 36644 45244 36650
rect 45192 36586 45244 36592
rect 44824 36236 44876 36242
rect 44824 36178 44876 36184
rect 44180 36032 44232 36038
rect 44180 35974 44232 35980
rect 43996 35692 44048 35698
rect 43996 35634 44048 35640
rect 43444 35624 43496 35630
rect 43444 35566 43496 35572
rect 43456 35290 43484 35566
rect 43444 35284 43496 35290
rect 43444 35226 43496 35232
rect 44008 34746 44036 35634
rect 43996 34740 44048 34746
rect 43996 34682 44048 34688
rect 44192 34610 44220 35974
rect 44836 35562 44864 36178
rect 44824 35556 44876 35562
rect 44824 35498 44876 35504
rect 44272 35080 44324 35086
rect 44272 35022 44324 35028
rect 44180 34604 44232 34610
rect 44180 34546 44232 34552
rect 43260 34060 43312 34066
rect 43260 34002 43312 34008
rect 43076 33992 43128 33998
rect 43076 33934 43128 33940
rect 43168 33992 43220 33998
rect 43168 33934 43220 33940
rect 42984 33516 43036 33522
rect 42984 33458 43036 33464
rect 42892 33108 42944 33114
rect 42892 33050 42944 33056
rect 42432 32904 42484 32910
rect 42432 32846 42484 32852
rect 42800 32904 42852 32910
rect 42800 32846 42852 32852
rect 42444 32434 42472 32846
rect 42616 32496 42668 32502
rect 42616 32438 42668 32444
rect 42432 32428 42484 32434
rect 42432 32370 42484 32376
rect 42064 32292 42116 32298
rect 42064 32234 42116 32240
rect 41328 32224 41380 32230
rect 41328 32166 41380 32172
rect 41340 31890 41368 32166
rect 42628 31958 42656 32438
rect 42708 32428 42760 32434
rect 42708 32370 42760 32376
rect 42616 31952 42668 31958
rect 42616 31894 42668 31900
rect 41328 31884 41380 31890
rect 41328 31826 41380 31832
rect 42628 31754 42656 31894
rect 41696 31748 41748 31754
rect 41696 31690 41748 31696
rect 42536 31726 42656 31754
rect 41708 31482 41736 31690
rect 41696 31476 41748 31482
rect 41696 31418 41748 31424
rect 42536 31346 42564 31726
rect 42524 31340 42576 31346
rect 42524 31282 42576 31288
rect 42720 30734 42748 32370
rect 42996 31346 43024 33458
rect 43088 32434 43116 33934
rect 43180 33658 43208 33934
rect 43168 33652 43220 33658
rect 43168 33594 43220 33600
rect 43076 32428 43128 32434
rect 43076 32370 43128 32376
rect 43272 31958 43300 34002
rect 43720 33856 43772 33862
rect 43720 33798 43772 33804
rect 43732 33590 43760 33798
rect 43720 33584 43772 33590
rect 43720 33526 43772 33532
rect 43628 33448 43680 33454
rect 43628 33390 43680 33396
rect 43640 33114 43668 33390
rect 43628 33108 43680 33114
rect 43628 33050 43680 33056
rect 44284 32910 44312 35022
rect 45204 33930 45232 36586
rect 45296 35086 45324 42570
rect 46296 41744 46348 41750
rect 46296 41686 46348 41692
rect 45376 41676 45428 41682
rect 45376 41618 45428 41624
rect 45388 41206 45416 41618
rect 45468 41608 45520 41614
rect 45468 41550 45520 41556
rect 45744 41608 45796 41614
rect 45744 41550 45796 41556
rect 45480 41460 45508 41550
rect 45652 41472 45704 41478
rect 45480 41432 45652 41460
rect 45652 41414 45704 41420
rect 45756 41274 45784 41550
rect 45744 41268 45796 41274
rect 45744 41210 45796 41216
rect 46308 41206 46336 41686
rect 46664 41540 46716 41546
rect 46664 41482 46716 41488
rect 45376 41200 45428 41206
rect 45376 41142 45428 41148
rect 46296 41200 46348 41206
rect 46296 41142 46348 41148
rect 45388 39914 45416 41142
rect 45928 41132 45980 41138
rect 45928 41074 45980 41080
rect 45940 41018 45968 41074
rect 46296 41064 46348 41070
rect 45940 41012 46296 41018
rect 45940 41006 46348 41012
rect 46386 41032 46442 41041
rect 45940 40990 46336 41006
rect 46386 40967 46388 40976
rect 46440 40967 46442 40976
rect 46388 40938 46440 40944
rect 45744 40928 45796 40934
rect 45744 40870 45796 40876
rect 45756 40526 45784 40870
rect 46676 40594 46704 41482
rect 47412 41414 47440 71318
rect 47646 71200 47758 71318
rect 48934 71200 49046 72000
rect 50222 71200 50334 72000
rect 51510 71200 51622 72000
rect 52798 71200 52910 72000
rect 54086 71346 54198 72000
rect 53852 71318 54198 71346
rect 48976 68898 49004 71200
rect 50264 69850 50292 71200
rect 50172 69822 50292 69850
rect 48976 68870 49280 68898
rect 48964 68808 49016 68814
rect 48964 68750 49016 68756
rect 48976 68338 49004 68750
rect 48964 68332 49016 68338
rect 48964 68274 49016 68280
rect 47584 56772 47636 56778
rect 47584 56714 47636 56720
rect 47596 55418 47624 56714
rect 48228 56704 48280 56710
rect 48228 56646 48280 56652
rect 48240 56370 48268 56646
rect 48228 56364 48280 56370
rect 48228 56306 48280 56312
rect 47768 56160 47820 56166
rect 47768 56102 47820 56108
rect 47584 55412 47636 55418
rect 47584 55354 47636 55360
rect 47780 55282 47808 56102
rect 48240 55826 48268 56306
rect 48780 56296 48832 56302
rect 48780 56238 48832 56244
rect 48792 55962 48820 56238
rect 48596 55956 48648 55962
rect 48596 55898 48648 55904
rect 48780 55956 48832 55962
rect 48780 55898 48832 55904
rect 48228 55820 48280 55826
rect 48228 55762 48280 55768
rect 48608 55758 48636 55898
rect 48596 55752 48648 55758
rect 48596 55694 48648 55700
rect 47952 55616 48004 55622
rect 47952 55558 48004 55564
rect 47768 55276 47820 55282
rect 47768 55218 47820 55224
rect 47676 54664 47728 54670
rect 47676 54606 47728 54612
rect 47688 54330 47716 54606
rect 47676 54324 47728 54330
rect 47676 54266 47728 54272
rect 47584 53780 47636 53786
rect 47584 53722 47636 53728
rect 47596 52494 47624 53722
rect 47964 53242 47992 55558
rect 48504 55276 48556 55282
rect 48504 55218 48556 55224
rect 48320 55072 48372 55078
rect 48320 55014 48372 55020
rect 48332 54670 48360 55014
rect 48320 54664 48372 54670
rect 48320 54606 48372 54612
rect 48516 54330 48544 55218
rect 48688 54528 48740 54534
rect 48688 54470 48740 54476
rect 48504 54324 48556 54330
rect 48504 54266 48556 54272
rect 48700 54194 48728 54470
rect 48688 54188 48740 54194
rect 48688 54130 48740 54136
rect 48700 53786 48728 54130
rect 48688 53780 48740 53786
rect 48688 53722 48740 53728
rect 48504 53576 48556 53582
rect 48504 53518 48556 53524
rect 48228 53508 48280 53514
rect 48228 53450 48280 53456
rect 47952 53236 48004 53242
rect 47952 53178 48004 53184
rect 48240 53106 48268 53450
rect 48516 53106 48544 53518
rect 48964 53440 49016 53446
rect 48964 53382 49016 53388
rect 47860 53100 47912 53106
rect 47860 53042 47912 53048
rect 48228 53100 48280 53106
rect 48228 53042 48280 53048
rect 48504 53100 48556 53106
rect 48504 53042 48556 53048
rect 47584 52488 47636 52494
rect 47584 52430 47636 52436
rect 47872 52426 47900 53042
rect 48228 52964 48280 52970
rect 48228 52906 48280 52912
rect 47860 52420 47912 52426
rect 47860 52362 47912 52368
rect 47584 52352 47636 52358
rect 47584 52294 47636 52300
rect 47596 52018 47624 52294
rect 47584 52012 47636 52018
rect 47584 51954 47636 51960
rect 48240 51814 48268 52906
rect 48976 52698 49004 53382
rect 48964 52692 49016 52698
rect 48964 52634 49016 52640
rect 48976 51882 49004 52634
rect 48964 51876 49016 51882
rect 48964 51818 49016 51824
rect 48228 51808 48280 51814
rect 48228 51750 48280 51756
rect 48240 50930 48268 51750
rect 48412 51400 48464 51406
rect 48412 51342 48464 51348
rect 47676 50924 47728 50930
rect 47676 50866 47728 50872
rect 48228 50924 48280 50930
rect 48228 50866 48280 50872
rect 47492 50176 47544 50182
rect 47492 50118 47544 50124
rect 47504 49366 47532 50118
rect 47688 49910 47716 50866
rect 48240 50386 48268 50866
rect 48424 50862 48452 51342
rect 48412 50856 48464 50862
rect 48412 50798 48464 50804
rect 48780 50856 48832 50862
rect 48780 50798 48832 50804
rect 48228 50380 48280 50386
rect 48228 50322 48280 50328
rect 47768 50312 47820 50318
rect 47768 50254 47820 50260
rect 47676 49904 47728 49910
rect 47596 49852 47676 49858
rect 47596 49846 47728 49852
rect 47596 49830 47716 49846
rect 47492 49360 47544 49366
rect 47492 49302 47544 49308
rect 47504 48006 47532 49302
rect 47596 48822 47624 49830
rect 47780 49774 47808 50254
rect 48320 50244 48372 50250
rect 48320 50186 48372 50192
rect 48136 50176 48188 50182
rect 48136 50118 48188 50124
rect 47768 49768 47820 49774
rect 47768 49710 47820 49716
rect 47676 49224 47728 49230
rect 47676 49166 47728 49172
rect 47688 48822 47716 49166
rect 48148 48890 48176 50118
rect 48228 49632 48280 49638
rect 48332 49586 48360 50186
rect 48280 49580 48360 49586
rect 48228 49574 48360 49580
rect 48240 49558 48360 49574
rect 48332 49434 48360 49558
rect 48320 49428 48372 49434
rect 48320 49370 48372 49376
rect 48136 48884 48188 48890
rect 48136 48826 48188 48832
rect 47584 48816 47636 48822
rect 47584 48758 47636 48764
rect 47676 48816 47728 48822
rect 47676 48758 47728 48764
rect 47596 48686 47624 48758
rect 47584 48680 47636 48686
rect 47584 48622 47636 48628
rect 47492 48000 47544 48006
rect 47492 47942 47544 47948
rect 47596 46714 47624 48622
rect 47952 48544 48004 48550
rect 47952 48486 48004 48492
rect 47964 48142 47992 48486
rect 47952 48136 48004 48142
rect 47952 48078 48004 48084
rect 47964 47734 47992 48078
rect 47952 47728 48004 47734
rect 47952 47670 48004 47676
rect 47584 46708 47636 46714
rect 47584 46650 47636 46656
rect 48044 46640 48096 46646
rect 48044 46582 48096 46588
rect 48056 45966 48084 46582
rect 48044 45960 48096 45966
rect 48044 45902 48096 45908
rect 47952 45484 48004 45490
rect 47952 45426 48004 45432
rect 47584 45280 47636 45286
rect 47584 45222 47636 45228
rect 47596 44946 47624 45222
rect 47584 44940 47636 44946
rect 47584 44882 47636 44888
rect 47676 44736 47728 44742
rect 47676 44678 47728 44684
rect 47688 44402 47716 44678
rect 47964 44538 47992 45426
rect 48056 45422 48084 45902
rect 48044 45416 48096 45422
rect 48044 45358 48096 45364
rect 48320 45280 48372 45286
rect 48320 45222 48372 45228
rect 48332 44878 48360 45222
rect 48320 44872 48372 44878
rect 48320 44814 48372 44820
rect 48424 44810 48452 50798
rect 48596 50720 48648 50726
rect 48596 50662 48648 50668
rect 48608 50318 48636 50662
rect 48792 50454 48820 50798
rect 49056 50720 49108 50726
rect 49056 50662 49108 50668
rect 49068 50522 49096 50662
rect 49056 50516 49108 50522
rect 49056 50458 49108 50464
rect 48780 50448 48832 50454
rect 48780 50390 48832 50396
rect 48596 50312 48648 50318
rect 48596 50254 48648 50260
rect 49068 49638 49096 50458
rect 49056 49632 49108 49638
rect 49056 49574 49108 49580
rect 48596 49224 48648 49230
rect 48596 49166 48648 49172
rect 48608 47666 48636 49166
rect 48688 48136 48740 48142
rect 48688 48078 48740 48084
rect 48700 47734 48728 48078
rect 49148 48068 49200 48074
rect 49148 48010 49200 48016
rect 49160 47734 49188 48010
rect 48688 47728 48740 47734
rect 48688 47670 48740 47676
rect 49148 47728 49200 47734
rect 49148 47670 49200 47676
rect 48596 47660 48648 47666
rect 48596 47602 48648 47608
rect 48504 45348 48556 45354
rect 48504 45290 48556 45296
rect 48412 44804 48464 44810
rect 48412 44746 48464 44752
rect 47952 44532 48004 44538
rect 47952 44474 48004 44480
rect 48516 44402 48544 45290
rect 47676 44396 47728 44402
rect 47676 44338 47728 44344
rect 47768 44396 47820 44402
rect 47768 44338 47820 44344
rect 48504 44396 48556 44402
rect 48504 44338 48556 44344
rect 48688 44396 48740 44402
rect 48688 44338 48740 44344
rect 47676 43648 47728 43654
rect 47676 43590 47728 43596
rect 47688 43314 47716 43590
rect 47780 43314 47808 44338
rect 48320 43716 48372 43722
rect 48320 43658 48372 43664
rect 47676 43308 47728 43314
rect 47676 43250 47728 43256
rect 47768 43308 47820 43314
rect 47768 43250 47820 43256
rect 48136 43104 48188 43110
rect 48136 43046 48188 43052
rect 48148 42702 48176 43046
rect 48136 42696 48188 42702
rect 48136 42638 48188 42644
rect 48332 42566 48360 43658
rect 48516 43450 48544 44338
rect 48596 44192 48648 44198
rect 48596 44134 48648 44140
rect 48608 43790 48636 44134
rect 48596 43784 48648 43790
rect 48596 43726 48648 43732
rect 48504 43444 48556 43450
rect 48504 43386 48556 43392
rect 48700 43314 48728 44338
rect 48688 43308 48740 43314
rect 48688 43250 48740 43256
rect 48320 42560 48372 42566
rect 48320 42502 48372 42508
rect 48596 42152 48648 42158
rect 48596 42094 48648 42100
rect 48608 41478 48636 42094
rect 48780 41608 48832 41614
rect 48780 41550 48832 41556
rect 48596 41472 48648 41478
rect 48596 41414 48648 41420
rect 47320 41386 47440 41414
rect 46664 40588 46716 40594
rect 46664 40530 46716 40536
rect 45744 40520 45796 40526
rect 45744 40462 45796 40468
rect 46112 40384 46164 40390
rect 46112 40326 46164 40332
rect 45376 39908 45428 39914
rect 45376 39850 45428 39856
rect 45388 39574 45416 39850
rect 45376 39568 45428 39574
rect 45376 39510 45428 39516
rect 45388 36922 45416 39510
rect 46124 39438 46152 40326
rect 46296 40180 46348 40186
rect 46296 40122 46348 40128
rect 46308 40050 46336 40122
rect 46296 40044 46348 40050
rect 46296 39986 46348 39992
rect 46572 40044 46624 40050
rect 46572 39986 46624 39992
rect 46584 39642 46612 39986
rect 46572 39636 46624 39642
rect 46572 39578 46624 39584
rect 46676 39506 46704 40530
rect 46756 40044 46808 40050
rect 46756 39986 46808 39992
rect 46664 39500 46716 39506
rect 46664 39442 46716 39448
rect 45652 39432 45704 39438
rect 45650 39400 45652 39409
rect 46112 39432 46164 39438
rect 45704 39400 45706 39409
rect 46112 39374 46164 39380
rect 45650 39335 45706 39344
rect 46020 39296 46072 39302
rect 46020 39238 46072 39244
rect 45836 39092 45888 39098
rect 45836 39034 45888 39040
rect 45848 38418 45876 39034
rect 46032 38418 46060 39238
rect 46676 39030 46704 39442
rect 46768 39409 46796 39986
rect 46848 39840 46900 39846
rect 46848 39782 46900 39788
rect 46860 39438 46888 39782
rect 46848 39432 46900 39438
rect 46754 39400 46810 39409
rect 46848 39374 46900 39380
rect 46754 39335 46810 39344
rect 46664 39024 46716 39030
rect 46664 38966 46716 38972
rect 45836 38412 45888 38418
rect 45836 38354 45888 38360
rect 46020 38412 46072 38418
rect 46020 38354 46072 38360
rect 46572 37800 46624 37806
rect 46572 37742 46624 37748
rect 46584 37126 46612 37742
rect 46572 37120 46624 37126
rect 46572 37062 46624 37068
rect 45376 36916 45428 36922
rect 45376 36858 45428 36864
rect 46768 36786 46796 39335
rect 47320 37942 47348 41386
rect 48044 41064 48096 41070
rect 48044 41006 48096 41012
rect 48056 40730 48084 41006
rect 48044 40724 48096 40730
rect 48044 40666 48096 40672
rect 48056 38962 48084 40666
rect 48792 40526 48820 41550
rect 48872 41472 48924 41478
rect 48872 41414 48924 41420
rect 48884 41206 48912 41414
rect 48872 41200 48924 41206
rect 48872 41142 48924 41148
rect 48780 40520 48832 40526
rect 48780 40462 48832 40468
rect 48136 40112 48188 40118
rect 48136 40054 48188 40060
rect 48148 39642 48176 40054
rect 48136 39636 48188 39642
rect 48136 39578 48188 39584
rect 48792 39438 48820 40462
rect 48964 40384 49016 40390
rect 48964 40326 49016 40332
rect 48976 40118 49004 40326
rect 48964 40112 49016 40118
rect 48964 40054 49016 40060
rect 48780 39432 48832 39438
rect 48780 39374 48832 39380
rect 48964 39296 49016 39302
rect 48964 39238 49016 39244
rect 48976 39030 49004 39238
rect 48964 39024 49016 39030
rect 48964 38966 49016 38972
rect 48044 38956 48096 38962
rect 48044 38898 48096 38904
rect 47584 38276 47636 38282
rect 47584 38218 47636 38224
rect 47308 37936 47360 37942
rect 47308 37878 47360 37884
rect 46848 37664 46900 37670
rect 46848 37606 46900 37612
rect 46860 37262 46888 37606
rect 46848 37256 46900 37262
rect 46848 37198 46900 37204
rect 45652 36780 45704 36786
rect 45652 36722 45704 36728
rect 46388 36780 46440 36786
rect 46388 36722 46440 36728
rect 46756 36780 46808 36786
rect 46756 36722 46808 36728
rect 45560 36168 45612 36174
rect 45560 36110 45612 36116
rect 45284 35080 45336 35086
rect 45284 35022 45336 35028
rect 45376 34740 45428 34746
rect 45376 34682 45428 34688
rect 45388 33998 45416 34682
rect 45572 34610 45600 36110
rect 45664 35222 45692 36722
rect 46400 36378 46428 36722
rect 46768 36650 46796 36722
rect 46756 36644 46808 36650
rect 46756 36586 46808 36592
rect 46572 36576 46624 36582
rect 46572 36518 46624 36524
rect 46388 36372 46440 36378
rect 46388 36314 46440 36320
rect 46584 36174 46612 36518
rect 46572 36168 46624 36174
rect 46572 36110 46624 36116
rect 46860 35698 46888 37198
rect 46848 35692 46900 35698
rect 46848 35634 46900 35640
rect 45652 35216 45704 35222
rect 46860 35170 46888 35634
rect 45652 35158 45704 35164
rect 45560 34604 45612 34610
rect 45560 34546 45612 34552
rect 45376 33992 45428 33998
rect 45376 33934 45428 33940
rect 44456 33924 44508 33930
rect 44456 33866 44508 33872
rect 45192 33924 45244 33930
rect 45192 33866 45244 33872
rect 43444 32904 43496 32910
rect 43444 32846 43496 32852
rect 44272 32904 44324 32910
rect 44272 32846 44324 32852
rect 43352 32224 43404 32230
rect 43352 32166 43404 32172
rect 43260 31952 43312 31958
rect 43260 31894 43312 31900
rect 42984 31340 43036 31346
rect 42984 31282 43036 31288
rect 42708 30728 42760 30734
rect 42708 30670 42760 30676
rect 41420 30592 41472 30598
rect 41420 30534 41472 30540
rect 42984 30592 43036 30598
rect 42984 30534 43036 30540
rect 41432 30326 41460 30534
rect 41420 30320 41472 30326
rect 41420 30262 41472 30268
rect 42996 30258 43024 30534
rect 43272 30326 43300 31894
rect 43364 31822 43392 32166
rect 43352 31816 43404 31822
rect 43352 31758 43404 31764
rect 43456 31686 43484 32846
rect 43720 32768 43772 32774
rect 43720 32710 43772 32716
rect 43732 32502 43760 32710
rect 44468 32586 44496 33866
rect 44468 32558 44680 32586
rect 43720 32496 43772 32502
rect 43720 32438 43772 32444
rect 43628 32428 43680 32434
rect 43628 32370 43680 32376
rect 43640 31890 43668 32370
rect 43628 31884 43680 31890
rect 43628 31826 43680 31832
rect 43444 31680 43496 31686
rect 43444 31622 43496 31628
rect 43456 31346 43484 31622
rect 43444 31340 43496 31346
rect 43444 31282 43496 31288
rect 43260 30320 43312 30326
rect 43260 30262 43312 30268
rect 42984 30252 43036 30258
rect 42984 30194 43036 30200
rect 43272 30138 43300 30262
rect 43640 30190 43668 31826
rect 43180 30110 43300 30138
rect 43628 30184 43680 30190
rect 43628 30126 43680 30132
rect 43180 29714 43208 30110
rect 43260 30048 43312 30054
rect 43260 29990 43312 29996
rect 43168 29708 43220 29714
rect 43168 29650 43220 29656
rect 43272 29170 43300 29990
rect 43640 29646 43668 30126
rect 43628 29640 43680 29646
rect 43628 29582 43680 29588
rect 43732 29170 43760 32438
rect 44364 32428 44416 32434
rect 44364 32370 44416 32376
rect 44376 32230 44404 32370
rect 44364 32224 44416 32230
rect 44364 32166 44416 32172
rect 44468 31754 44496 32558
rect 44548 32428 44600 32434
rect 44548 32370 44600 32376
rect 44560 32026 44588 32370
rect 44652 32366 44680 32558
rect 45572 32502 45600 34546
rect 45664 33998 45692 35158
rect 46768 35142 46888 35170
rect 46768 34610 46796 35142
rect 47492 35080 47544 35086
rect 47492 35022 47544 35028
rect 47504 34746 47532 35022
rect 47492 34740 47544 34746
rect 47492 34682 47544 34688
rect 45744 34604 45796 34610
rect 45744 34546 45796 34552
rect 46756 34604 46808 34610
rect 46756 34546 46808 34552
rect 45756 34202 45784 34546
rect 45744 34196 45796 34202
rect 45744 34138 45796 34144
rect 45652 33992 45704 33998
rect 45652 33934 45704 33940
rect 46768 33522 46796 34546
rect 46756 33516 46808 33522
rect 46756 33458 46808 33464
rect 46768 33402 46796 33458
rect 46768 33374 46888 33402
rect 46756 32904 46808 32910
rect 46756 32846 46808 32852
rect 45560 32496 45612 32502
rect 45560 32438 45612 32444
rect 44640 32360 44692 32366
rect 44640 32302 44692 32308
rect 46768 32230 46796 32846
rect 46756 32224 46808 32230
rect 46756 32166 46808 32172
rect 44548 32020 44600 32026
rect 44548 31962 44600 31968
rect 44376 31726 44496 31754
rect 44180 31340 44232 31346
rect 44180 31282 44232 31288
rect 43996 31272 44048 31278
rect 43996 31214 44048 31220
rect 43904 31136 43956 31142
rect 43904 31078 43956 31084
rect 43916 30258 43944 31078
rect 44008 30734 44036 31214
rect 44192 30938 44220 31282
rect 44180 30932 44232 30938
rect 44180 30874 44232 30880
rect 43996 30728 44048 30734
rect 43996 30670 44048 30676
rect 43904 30252 43956 30258
rect 43904 30194 43956 30200
rect 44272 29504 44324 29510
rect 44272 29446 44324 29452
rect 44284 29238 44312 29446
rect 44376 29306 44404 31726
rect 44456 31136 44508 31142
rect 44456 31078 44508 31084
rect 44468 30326 44496 31078
rect 45468 30660 45520 30666
rect 45468 30602 45520 30608
rect 45480 30394 45508 30602
rect 45468 30388 45520 30394
rect 45468 30330 45520 30336
rect 44456 30320 44508 30326
rect 44456 30262 44508 30268
rect 46860 29646 46888 33374
rect 46940 33312 46992 33318
rect 46940 33254 46992 33260
rect 46952 32978 46980 33254
rect 46940 32972 46992 32978
rect 46940 32914 46992 32920
rect 47596 31754 47624 38218
rect 48044 37936 48096 37942
rect 48044 37878 48096 37884
rect 48056 37806 48084 37878
rect 47768 37800 47820 37806
rect 47768 37742 47820 37748
rect 48044 37800 48096 37806
rect 48044 37742 48096 37748
rect 47780 37466 47808 37742
rect 47768 37460 47820 37466
rect 47768 37402 47820 37408
rect 47860 36712 47912 36718
rect 47860 36654 47912 36660
rect 47872 36378 47900 36654
rect 47860 36372 47912 36378
rect 47860 36314 47912 36320
rect 47872 35698 47900 36314
rect 47860 35692 47912 35698
rect 47860 35634 47912 35640
rect 49252 35154 49280 68870
rect 50172 68202 50200 69822
rect 50294 69660 50602 69680
rect 50294 69658 50300 69660
rect 50356 69658 50380 69660
rect 50436 69658 50460 69660
rect 50516 69658 50540 69660
rect 50596 69658 50602 69660
rect 50356 69606 50358 69658
rect 50538 69606 50540 69658
rect 50294 69604 50300 69606
rect 50356 69604 50380 69606
rect 50436 69604 50460 69606
rect 50516 69604 50540 69606
rect 50596 69604 50602 69606
rect 50294 69584 50602 69604
rect 50712 69216 50764 69222
rect 50712 69158 50764 69164
rect 50724 68882 50752 69158
rect 51552 68882 51580 71200
rect 52840 68950 52868 71200
rect 52920 69216 52972 69222
rect 52920 69158 52972 69164
rect 52828 68944 52880 68950
rect 52828 68886 52880 68892
rect 52932 68882 52960 69158
rect 50712 68876 50764 68882
rect 50712 68818 50764 68824
rect 51540 68876 51592 68882
rect 51540 68818 51592 68824
rect 52920 68876 52972 68882
rect 52920 68818 52972 68824
rect 52920 68740 52972 68746
rect 52920 68682 52972 68688
rect 50294 68572 50602 68592
rect 50294 68570 50300 68572
rect 50356 68570 50380 68572
rect 50436 68570 50460 68572
rect 50516 68570 50540 68572
rect 50596 68570 50602 68572
rect 50356 68518 50358 68570
rect 50538 68518 50540 68570
rect 50294 68516 50300 68518
rect 50356 68516 50380 68518
rect 50436 68516 50460 68518
rect 50516 68516 50540 68518
rect 50596 68516 50602 68518
rect 50294 68496 50602 68516
rect 52932 68474 52960 68682
rect 52920 68468 52972 68474
rect 52920 68410 52972 68416
rect 52736 68332 52788 68338
rect 52736 68274 52788 68280
rect 50252 68264 50304 68270
rect 50252 68206 50304 68212
rect 50160 68196 50212 68202
rect 50160 68138 50212 68144
rect 50264 67930 50292 68206
rect 50252 67924 50304 67930
rect 50252 67866 50304 67872
rect 50160 67720 50212 67726
rect 50160 67662 50212 67668
rect 50172 66638 50200 67662
rect 50294 67484 50602 67504
rect 50294 67482 50300 67484
rect 50356 67482 50380 67484
rect 50436 67482 50460 67484
rect 50516 67482 50540 67484
rect 50596 67482 50602 67484
rect 50356 67430 50358 67482
rect 50538 67430 50540 67482
rect 50294 67428 50300 67430
rect 50356 67428 50380 67430
rect 50436 67428 50460 67430
rect 50516 67428 50540 67430
rect 50596 67428 50602 67430
rect 50294 67408 50602 67428
rect 50160 66632 50212 66638
rect 50160 66574 50212 66580
rect 50172 65210 50200 66574
rect 50294 66396 50602 66416
rect 50294 66394 50300 66396
rect 50356 66394 50380 66396
rect 50436 66394 50460 66396
rect 50516 66394 50540 66396
rect 50596 66394 50602 66396
rect 50356 66342 50358 66394
rect 50538 66342 50540 66394
rect 50294 66340 50300 66342
rect 50356 66340 50380 66342
rect 50436 66340 50460 66342
rect 50516 66340 50540 66342
rect 50596 66340 50602 66342
rect 50294 66320 50602 66340
rect 52748 66162 52776 68274
rect 52736 66156 52788 66162
rect 52736 66098 52788 66104
rect 53104 66156 53156 66162
rect 53104 66098 53156 66104
rect 50294 65308 50602 65328
rect 50294 65306 50300 65308
rect 50356 65306 50380 65308
rect 50436 65306 50460 65308
rect 50516 65306 50540 65308
rect 50596 65306 50602 65308
rect 50356 65254 50358 65306
rect 50538 65254 50540 65306
rect 50294 65252 50300 65254
rect 50356 65252 50380 65254
rect 50436 65252 50460 65254
rect 50516 65252 50540 65254
rect 50596 65252 50602 65254
rect 50294 65232 50602 65252
rect 50160 65204 50212 65210
rect 50160 65146 50212 65152
rect 50294 64220 50602 64240
rect 50294 64218 50300 64220
rect 50356 64218 50380 64220
rect 50436 64218 50460 64220
rect 50516 64218 50540 64220
rect 50596 64218 50602 64220
rect 50356 64166 50358 64218
rect 50538 64166 50540 64218
rect 50294 64164 50300 64166
rect 50356 64164 50380 64166
rect 50436 64164 50460 64166
rect 50516 64164 50540 64166
rect 50596 64164 50602 64166
rect 50294 64144 50602 64164
rect 50294 63132 50602 63152
rect 50294 63130 50300 63132
rect 50356 63130 50380 63132
rect 50436 63130 50460 63132
rect 50516 63130 50540 63132
rect 50596 63130 50602 63132
rect 50356 63078 50358 63130
rect 50538 63078 50540 63130
rect 50294 63076 50300 63078
rect 50356 63076 50380 63078
rect 50436 63076 50460 63078
rect 50516 63076 50540 63078
rect 50596 63076 50602 63078
rect 50294 63056 50602 63076
rect 50294 62044 50602 62064
rect 50294 62042 50300 62044
rect 50356 62042 50380 62044
rect 50436 62042 50460 62044
rect 50516 62042 50540 62044
rect 50596 62042 50602 62044
rect 50356 61990 50358 62042
rect 50538 61990 50540 62042
rect 50294 61988 50300 61990
rect 50356 61988 50380 61990
rect 50436 61988 50460 61990
rect 50516 61988 50540 61990
rect 50596 61988 50602 61990
rect 50294 61968 50602 61988
rect 50294 60956 50602 60976
rect 50294 60954 50300 60956
rect 50356 60954 50380 60956
rect 50436 60954 50460 60956
rect 50516 60954 50540 60956
rect 50596 60954 50602 60956
rect 50356 60902 50358 60954
rect 50538 60902 50540 60954
rect 50294 60900 50300 60902
rect 50356 60900 50380 60902
rect 50436 60900 50460 60902
rect 50516 60900 50540 60902
rect 50596 60900 50602 60902
rect 50294 60880 50602 60900
rect 50294 59868 50602 59888
rect 50294 59866 50300 59868
rect 50356 59866 50380 59868
rect 50436 59866 50460 59868
rect 50516 59866 50540 59868
rect 50596 59866 50602 59868
rect 50356 59814 50358 59866
rect 50538 59814 50540 59866
rect 50294 59812 50300 59814
rect 50356 59812 50380 59814
rect 50436 59812 50460 59814
rect 50516 59812 50540 59814
rect 50596 59812 50602 59814
rect 50294 59792 50602 59812
rect 50294 58780 50602 58800
rect 50294 58778 50300 58780
rect 50356 58778 50380 58780
rect 50436 58778 50460 58780
rect 50516 58778 50540 58780
rect 50596 58778 50602 58780
rect 50356 58726 50358 58778
rect 50538 58726 50540 58778
rect 50294 58724 50300 58726
rect 50356 58724 50380 58726
rect 50436 58724 50460 58726
rect 50516 58724 50540 58726
rect 50596 58724 50602 58726
rect 50294 58704 50602 58724
rect 50294 57692 50602 57712
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57616 50602 57636
rect 53116 57458 53144 66098
rect 53852 59702 53880 71318
rect 54086 71200 54198 71318
rect 55374 71200 55486 72000
rect 56662 71200 56774 72000
rect 57950 71200 58062 72000
rect 59238 71200 59350 72000
rect 60526 71200 60638 72000
rect 61814 71346 61926 72000
rect 60752 71318 61926 71346
rect 55416 69426 55444 71200
rect 55404 69420 55456 69426
rect 55404 69362 55456 69368
rect 55680 69216 55732 69222
rect 55680 69158 55732 69164
rect 56508 69216 56560 69222
rect 56508 69158 56560 69164
rect 53840 59696 53892 59702
rect 53840 59638 53892 59644
rect 53104 57452 53156 57458
rect 53104 57394 53156 57400
rect 50620 56840 50672 56846
rect 50620 56782 50672 56788
rect 50160 56704 50212 56710
rect 50160 56646 50212 56652
rect 50172 56438 50200 56646
rect 50294 56604 50602 56624
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56528 50602 56548
rect 50160 56432 50212 56438
rect 50160 56374 50212 56380
rect 49700 56364 49752 56370
rect 49700 56306 49752 56312
rect 50344 56364 50396 56370
rect 50344 56306 50396 56312
rect 49712 54194 49740 56306
rect 50356 55758 50384 56306
rect 50528 56160 50580 56166
rect 50528 56102 50580 56108
rect 50540 55826 50568 56102
rect 50632 55962 50660 56782
rect 50620 55956 50672 55962
rect 50620 55898 50672 55904
rect 55692 55894 55720 69158
rect 56520 68882 56548 69158
rect 56704 68882 56732 71200
rect 57244 69420 57296 69426
rect 57244 69362 57296 69368
rect 56508 68876 56560 68882
rect 56508 68818 56560 68824
rect 56692 68876 56744 68882
rect 56692 68818 56744 68824
rect 56416 68740 56468 68746
rect 56416 68682 56468 68688
rect 56428 68474 56456 68682
rect 56416 68468 56468 68474
rect 56416 68410 56468 68416
rect 57256 68406 57284 69362
rect 57336 69216 57388 69222
rect 57336 69158 57388 69164
rect 57244 68400 57296 68406
rect 57244 68342 57296 68348
rect 56232 68332 56284 68338
rect 56232 68274 56284 68280
rect 56244 63034 56272 68274
rect 56232 63028 56284 63034
rect 56232 62970 56284 62976
rect 57256 62898 57284 68342
rect 57348 68338 57376 69158
rect 57336 68332 57388 68338
rect 57336 68274 57388 68280
rect 57992 68252 58020 71200
rect 59728 69352 59780 69358
rect 59728 69294 59780 69300
rect 58072 69216 58124 69222
rect 58072 69158 58124 69164
rect 58084 68406 58112 69158
rect 59740 68814 59768 69294
rect 60568 68950 60596 71200
rect 60648 69216 60700 69222
rect 60648 69158 60700 69164
rect 60556 68944 60608 68950
rect 60556 68886 60608 68892
rect 60660 68882 60688 69158
rect 60648 68876 60700 68882
rect 60648 68818 60700 68824
rect 59728 68808 59780 68814
rect 59728 68750 59780 68756
rect 59740 68678 59768 68750
rect 59728 68672 59780 68678
rect 59728 68614 59780 68620
rect 58072 68400 58124 68406
rect 58072 68342 58124 68348
rect 58072 68264 58124 68270
rect 57992 68224 58072 68252
rect 58072 68206 58124 68212
rect 57244 62892 57296 62898
rect 57244 62834 57296 62840
rect 55680 55888 55732 55894
rect 55680 55830 55732 55836
rect 50528 55820 50580 55826
rect 50528 55762 50580 55768
rect 50344 55752 50396 55758
rect 50344 55694 50396 55700
rect 50294 55516 50602 55536
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55440 50602 55460
rect 51264 55276 51316 55282
rect 51264 55218 51316 55224
rect 50436 55072 50488 55078
rect 50436 55014 50488 55020
rect 51080 55072 51132 55078
rect 51080 55014 51132 55020
rect 50448 54738 50476 55014
rect 50436 54732 50488 54738
rect 50436 54674 50488 54680
rect 51092 54670 51120 55014
rect 51080 54664 51132 54670
rect 51080 54606 51132 54612
rect 49884 54528 49936 54534
rect 49884 54470 49936 54476
rect 49700 54188 49752 54194
rect 49700 54130 49752 54136
rect 49896 54126 49924 54470
rect 50294 54428 50602 54448
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54352 50602 54372
rect 51276 54330 51304 55218
rect 51264 54324 51316 54330
rect 51264 54266 51316 54272
rect 50068 54188 50120 54194
rect 50068 54130 50120 54136
rect 50160 54188 50212 54194
rect 50160 54130 50212 54136
rect 49884 54120 49936 54126
rect 49884 54062 49936 54068
rect 49896 53718 49924 54062
rect 49884 53712 49936 53718
rect 49884 53654 49936 53660
rect 49884 53440 49936 53446
rect 49884 53382 49936 53388
rect 49896 53106 49924 53382
rect 50080 53106 50108 54130
rect 50172 53242 50200 54130
rect 50804 53984 50856 53990
rect 50804 53926 50856 53932
rect 50816 53582 50844 53926
rect 50620 53576 50672 53582
rect 50620 53518 50672 53524
rect 50804 53576 50856 53582
rect 50804 53518 50856 53524
rect 50294 53340 50602 53360
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53264 50602 53284
rect 50632 53242 50660 53518
rect 50160 53236 50212 53242
rect 50160 53178 50212 53184
rect 50620 53236 50672 53242
rect 50620 53178 50672 53184
rect 49884 53100 49936 53106
rect 49884 53042 49936 53048
rect 50068 53100 50120 53106
rect 50068 53042 50120 53048
rect 50712 53100 50764 53106
rect 50712 53042 50764 53048
rect 49792 52352 49844 52358
rect 49792 52294 49844 52300
rect 49804 52018 49832 52294
rect 49792 52012 49844 52018
rect 49792 51954 49844 51960
rect 50080 51474 50108 53042
rect 50724 52494 50752 53042
rect 50712 52488 50764 52494
rect 50712 52430 50764 52436
rect 50294 52252 50602 52272
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52176 50602 52196
rect 51080 52012 51132 52018
rect 51080 51954 51132 51960
rect 50528 51808 50580 51814
rect 50528 51750 50580 51756
rect 50540 51474 50568 51750
rect 51092 51542 51120 51954
rect 51080 51536 51132 51542
rect 51080 51478 51132 51484
rect 50068 51468 50120 51474
rect 50068 51410 50120 51416
rect 50528 51468 50580 51474
rect 50528 51410 50580 51416
rect 50540 51354 50568 51410
rect 50160 51332 50212 51338
rect 50540 51326 50660 51354
rect 50160 51274 50212 51280
rect 50172 50930 50200 51274
rect 50294 51164 50602 51184
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51088 50602 51108
rect 50160 50924 50212 50930
rect 50160 50866 50212 50872
rect 50068 50516 50120 50522
rect 50068 50458 50120 50464
rect 49792 50244 49844 50250
rect 49792 50186 49844 50192
rect 49332 49972 49384 49978
rect 49332 49914 49384 49920
rect 49344 49842 49372 49914
rect 49332 49836 49384 49842
rect 49332 49778 49384 49784
rect 49344 49230 49372 49778
rect 49332 49224 49384 49230
rect 49332 49166 49384 49172
rect 49424 48544 49476 48550
rect 49424 48486 49476 48492
rect 49700 48544 49752 48550
rect 49700 48486 49752 48492
rect 49436 48142 49464 48486
rect 49712 48210 49740 48486
rect 49700 48204 49752 48210
rect 49700 48146 49752 48152
rect 49424 48136 49476 48142
rect 49424 48078 49476 48084
rect 49700 47728 49752 47734
rect 49700 47670 49752 47676
rect 49712 46646 49740 47670
rect 49804 47598 49832 50186
rect 50080 49638 50108 50458
rect 50632 50318 50660 51326
rect 51540 50924 51592 50930
rect 51540 50866 51592 50872
rect 50988 50856 51040 50862
rect 50988 50798 51040 50804
rect 51000 50522 51028 50798
rect 50988 50516 51040 50522
rect 50988 50458 51040 50464
rect 50160 50312 50212 50318
rect 50160 50254 50212 50260
rect 50620 50312 50672 50318
rect 50620 50254 50672 50260
rect 51356 50312 51408 50318
rect 51356 50254 51408 50260
rect 50172 49960 50200 50254
rect 50294 50076 50602 50096
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50000 50602 50020
rect 50172 49932 50292 49960
rect 50264 49774 50292 49932
rect 50632 49842 50660 50254
rect 51368 49978 51396 50254
rect 51356 49972 51408 49978
rect 51356 49914 51408 49920
rect 50620 49836 50672 49842
rect 50620 49778 50672 49784
rect 51356 49836 51408 49842
rect 51356 49778 51408 49784
rect 50252 49768 50304 49774
rect 50252 49710 50304 49716
rect 50068 49632 50120 49638
rect 50068 49574 50120 49580
rect 50264 49230 50292 49710
rect 50252 49224 50304 49230
rect 50252 49166 50304 49172
rect 50294 48988 50602 49008
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48912 50602 48932
rect 51368 48754 51396 49778
rect 51552 49230 51580 50866
rect 52736 50720 52788 50726
rect 52736 50662 52788 50668
rect 52748 50318 52776 50662
rect 52736 50312 52788 50318
rect 52736 50254 52788 50260
rect 52092 49836 52144 49842
rect 52092 49778 52144 49784
rect 52000 49632 52052 49638
rect 52000 49574 52052 49580
rect 52012 49230 52040 49574
rect 52104 49434 52132 49778
rect 52092 49428 52144 49434
rect 52092 49370 52144 49376
rect 51540 49224 51592 49230
rect 51540 49166 51592 49172
rect 51632 49224 51684 49230
rect 51632 49166 51684 49172
rect 52000 49224 52052 49230
rect 52000 49166 52052 49172
rect 50160 48748 50212 48754
rect 50160 48690 50212 48696
rect 51356 48748 51408 48754
rect 51356 48690 51408 48696
rect 50172 48006 50200 48690
rect 50160 48000 50212 48006
rect 50160 47942 50212 47948
rect 50172 47734 50200 47942
rect 50294 47900 50602 47920
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47824 50602 47844
rect 50160 47728 50212 47734
rect 50160 47670 50212 47676
rect 50620 47660 50672 47666
rect 50620 47602 50672 47608
rect 49792 47592 49844 47598
rect 49792 47534 49844 47540
rect 50294 46812 50602 46832
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46736 50602 46756
rect 49700 46640 49752 46646
rect 49700 46582 49752 46588
rect 49424 46504 49476 46510
rect 49424 46446 49476 46452
rect 49436 46170 49464 46446
rect 49424 46164 49476 46170
rect 49424 46106 49476 46112
rect 50632 46034 50660 47602
rect 50804 47592 50856 47598
rect 50804 47534 50856 47540
rect 50816 46714 50844 47534
rect 51368 46986 51396 48690
rect 51448 47660 51500 47666
rect 51448 47602 51500 47608
rect 51460 47258 51488 47602
rect 51448 47252 51500 47258
rect 51448 47194 51500 47200
rect 51356 46980 51408 46986
rect 51356 46922 51408 46928
rect 50804 46708 50856 46714
rect 50804 46650 50856 46656
rect 50620 46028 50672 46034
rect 50620 45970 50672 45976
rect 50294 45724 50602 45744
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45648 50602 45668
rect 50160 45416 50212 45422
rect 50160 45358 50212 45364
rect 50632 45370 50660 45970
rect 50172 45082 50200 45358
rect 50632 45342 50844 45370
rect 50816 45286 50844 45342
rect 50804 45280 50856 45286
rect 50804 45222 50856 45228
rect 50160 45076 50212 45082
rect 50160 45018 50212 45024
rect 51368 44878 51396 46922
rect 51460 46578 51488 47194
rect 51552 46594 51580 49166
rect 51644 48890 51672 49166
rect 51632 48884 51684 48890
rect 51632 48826 51684 48832
rect 51632 47660 51684 47666
rect 51632 47602 51684 47608
rect 51644 46714 51672 47602
rect 51724 47456 51776 47462
rect 51724 47398 51776 47404
rect 51736 47054 51764 47398
rect 51724 47048 51776 47054
rect 51724 46990 51776 46996
rect 58716 46980 58768 46986
rect 58716 46922 58768 46928
rect 51632 46708 51684 46714
rect 51632 46650 51684 46656
rect 51552 46578 51764 46594
rect 51448 46572 51500 46578
rect 51552 46572 51776 46578
rect 51552 46566 51724 46572
rect 51448 46514 51500 46520
rect 51724 46514 51776 46520
rect 51736 45898 51764 46514
rect 51724 45892 51776 45898
rect 51724 45834 51776 45840
rect 51448 45824 51500 45830
rect 51448 45766 51500 45772
rect 51460 45558 51488 45766
rect 51448 45552 51500 45558
rect 51448 45494 51500 45500
rect 51356 44872 51408 44878
rect 51356 44814 51408 44820
rect 50294 44636 50602 44656
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44560 50602 44580
rect 51368 44538 51396 44814
rect 51356 44532 51408 44538
rect 51356 44474 51408 44480
rect 50294 43548 50602 43568
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43472 50602 43492
rect 50294 42460 50602 42480
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42384 50602 42404
rect 49424 42152 49476 42158
rect 49424 42094 49476 42100
rect 49436 41750 49464 42094
rect 58728 41818 58756 46922
rect 58716 41812 58768 41818
rect 58716 41754 58768 41760
rect 49424 41744 49476 41750
rect 49424 41686 49476 41692
rect 50294 41372 50602 41392
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41296 50602 41316
rect 50294 40284 50602 40304
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40208 50602 40228
rect 50294 39196 50602 39216
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39120 50602 39140
rect 50620 38888 50672 38894
rect 50620 38830 50672 38836
rect 50068 38208 50120 38214
rect 50068 38150 50120 38156
rect 50080 37942 50108 38150
rect 50294 38108 50602 38128
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38032 50602 38052
rect 50068 37936 50120 37942
rect 50068 37878 50120 37884
rect 50294 37020 50602 37040
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36944 50602 36964
rect 50294 35932 50602 35952
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35856 50602 35876
rect 49608 35624 49660 35630
rect 49608 35566 49660 35572
rect 49240 35148 49292 35154
rect 49240 35090 49292 35096
rect 47676 35012 47728 35018
rect 47676 34954 47728 34960
rect 47688 34746 47716 34954
rect 47676 34740 47728 34746
rect 47676 34682 47728 34688
rect 47596 31726 47716 31754
rect 46848 29640 46900 29646
rect 46848 29582 46900 29588
rect 44364 29300 44416 29306
rect 44364 29242 44416 29248
rect 44272 29232 44324 29238
rect 44272 29174 44324 29180
rect 43260 29164 43312 29170
rect 43260 29106 43312 29112
rect 43720 29164 43772 29170
rect 43720 29106 43772 29112
rect 43732 29034 43760 29106
rect 41512 29028 41564 29034
rect 41512 28970 41564 28976
rect 43720 29028 43772 29034
rect 43720 28970 43772 28976
rect 44180 29028 44232 29034
rect 44180 28970 44232 28976
rect 41524 28082 41552 28970
rect 42892 28960 42944 28966
rect 42892 28902 42944 28908
rect 42904 28558 42932 28902
rect 44192 28762 44220 28970
rect 44180 28756 44232 28762
rect 44180 28698 44232 28704
rect 42892 28552 42944 28558
rect 42892 28494 42944 28500
rect 44376 28150 44404 29242
rect 45928 29096 45980 29102
rect 45928 29038 45980 29044
rect 44364 28144 44416 28150
rect 44364 28086 44416 28092
rect 41512 28076 41564 28082
rect 41512 28018 41564 28024
rect 41512 27328 41564 27334
rect 41512 27270 41564 27276
rect 41524 26450 41552 27270
rect 45744 26784 45796 26790
rect 45744 26726 45796 26732
rect 40868 26444 40920 26450
rect 40868 26386 40920 26392
rect 41236 26444 41288 26450
rect 41236 26386 41288 26392
rect 41512 26444 41564 26450
rect 41512 26386 41564 26392
rect 43168 26308 43220 26314
rect 43168 26250 43220 26256
rect 43180 16590 43208 26250
rect 43168 16584 43220 16590
rect 38856 16546 39528 16574
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34612 4140 34664 4146
rect 34612 4082 34664 4088
rect 36084 4140 36136 4146
rect 36084 4082 36136 4088
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 33416 3052 33468 3058
rect 33416 2994 33468 3000
rect 32312 2644 32364 2650
rect 32312 2586 32364 2592
rect 33428 2514 33456 2994
rect 34612 2984 34664 2990
rect 34612 2926 34664 2932
rect 34796 2984 34848 2990
rect 34796 2926 34848 2932
rect 34624 2650 34652 2926
rect 34612 2644 34664 2650
rect 34612 2586 34664 2592
rect 33416 2508 33468 2514
rect 33416 2450 33468 2456
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 32128 2304 32180 2310
rect 32128 2246 32180 2252
rect 32232 800 32260 2382
rect 34808 800 34836 2926
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 36096 800 36124 4082
rect 38108 3528 38160 3534
rect 38108 3470 38160 3476
rect 37280 3188 37332 3194
rect 37280 3130 37332 3136
rect 37292 2446 37320 3130
rect 38120 3058 38148 3470
rect 38108 3052 38160 3058
rect 38108 2994 38160 3000
rect 38292 2984 38344 2990
rect 38292 2926 38344 2932
rect 38660 2984 38712 2990
rect 38660 2926 38712 2932
rect 38304 2650 38332 2926
rect 38292 2644 38344 2650
rect 38292 2586 38344 2592
rect 37280 2440 37332 2446
rect 37280 2382 37332 2388
rect 38672 800 38700 2926
rect 2870 776 2926 785
rect 2870 711 2926 720
rect 3210 0 3322 800
rect 4498 0 4610 800
rect 5786 0 5898 800
rect 7074 0 7186 800
rect 8362 0 8474 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 12226 0 12338 800
rect 13514 0 13626 800
rect 14802 0 14914 800
rect 16090 0 16202 800
rect 17378 0 17490 800
rect 18666 0 18778 800
rect 19954 0 20066 800
rect 21242 0 21354 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 24462 0 24574 800
rect 25750 0 25862 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 29614 0 29726 800
rect 30902 0 31014 800
rect 32190 0 32302 800
rect 33478 0 33590 800
rect 34766 0 34878 800
rect 36054 0 36166 800
rect 37342 0 37454 800
rect 38630 0 38742 800
rect 39500 762 39528 16546
rect 43168 16526 43220 16532
rect 45756 4146 45784 26726
rect 45744 4140 45796 4146
rect 45744 4082 45796 4088
rect 45940 4078 45968 29038
rect 41236 4072 41288 4078
rect 41236 4014 41288 4020
rect 45928 4072 45980 4078
rect 45928 4014 45980 4020
rect 39776 870 39988 898
rect 39776 762 39804 870
rect 39960 800 39988 870
rect 41248 800 41276 4014
rect 46388 3936 46440 3942
rect 46388 3878 46440 3884
rect 46400 3602 46428 3878
rect 47688 3670 47716 31726
rect 49620 30326 49648 35566
rect 50294 34844 50602 34864
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34768 50602 34788
rect 50294 33756 50602 33776
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33680 50602 33700
rect 50294 32668 50602 32688
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32592 50602 32612
rect 50294 31580 50602 31600
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31504 50602 31524
rect 50294 30492 50602 30512
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30416 50602 30436
rect 49608 30320 49660 30326
rect 49608 30262 49660 30268
rect 50294 29404 50602 29424
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29328 50602 29348
rect 50294 28316 50602 28336
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28240 50602 28260
rect 50294 27228 50602 27248
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27152 50602 27172
rect 50294 26140 50602 26160
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26064 50602 26084
rect 50294 25052 50602 25072
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24976 50602 24996
rect 50294 23964 50602 23984
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23888 50602 23908
rect 50294 22876 50602 22896
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22800 50602 22820
rect 50294 21788 50602 21808
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21712 50602 21732
rect 50294 20700 50602 20720
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20624 50602 20644
rect 50294 19612 50602 19632
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19536 50602 19556
rect 50294 18524 50602 18544
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18448 50602 18468
rect 50294 17436 50602 17456
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17360 50602 17380
rect 50294 16348 50602 16368
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16272 50602 16292
rect 50294 15260 50602 15280
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15184 50602 15204
rect 50294 14172 50602 14192
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14096 50602 14116
rect 50294 13084 50602 13104
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13008 50602 13028
rect 50294 11996 50602 12016
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11920 50602 11940
rect 50294 10908 50602 10928
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10832 50602 10852
rect 50294 9820 50602 9840
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9744 50602 9764
rect 50294 8732 50602 8752
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8656 50602 8676
rect 50294 7644 50602 7664
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7568 50602 7588
rect 50294 6556 50602 6576
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6480 50602 6500
rect 50294 5468 50602 5488
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5392 50602 5412
rect 50294 4380 50602 4400
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4304 50602 4324
rect 47676 3664 47728 3670
rect 47676 3606 47728 3612
rect 46388 3596 46440 3602
rect 46388 3538 46440 3544
rect 47032 3596 47084 3602
rect 47032 3538 47084 3544
rect 46204 3528 46256 3534
rect 46204 3470 46256 3476
rect 43812 3460 43864 3466
rect 43812 3402 43864 3408
rect 42524 2372 42576 2378
rect 42524 2314 42576 2320
rect 42536 800 42564 2314
rect 43824 800 43852 3402
rect 44824 3392 44876 3398
rect 44824 3334 44876 3340
rect 44836 3126 44864 3334
rect 44824 3120 44876 3126
rect 44824 3062 44876 3068
rect 45100 2984 45152 2990
rect 45100 2926 45152 2932
rect 45112 800 45140 2926
rect 46216 2650 46244 3470
rect 46204 2644 46256 2650
rect 46204 2586 46256 2592
rect 47044 800 47072 3538
rect 50294 3292 50602 3312
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3216 50602 3236
rect 50294 2204 50602 2224
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2128 50602 2148
rect 50632 1358 50660 38830
rect 51724 37800 51776 37806
rect 51724 37742 51776 37748
rect 51736 3534 51764 37742
rect 59740 3534 59768 68614
rect 60752 41070 60780 71318
rect 61814 71200 61926 71318
rect 63102 71200 63214 72000
rect 64390 71200 64502 72000
rect 65678 71200 65790 72000
rect 66966 71200 67078 72000
rect 68254 71200 68366 72000
rect 69542 71200 69654 72000
rect 62212 69216 62264 69222
rect 62212 69158 62264 69164
rect 62224 68882 62252 69158
rect 63144 68882 63172 71200
rect 65720 69442 65748 71200
rect 64892 69414 65748 69442
rect 62212 68876 62264 68882
rect 62212 68818 62264 68824
rect 63132 68876 63184 68882
rect 63132 68818 63184 68824
rect 62948 68740 63000 68746
rect 62948 68682 63000 68688
rect 62960 68474 62988 68682
rect 62948 68468 63000 68474
rect 62948 68410 63000 68416
rect 61568 68332 61620 68338
rect 61568 68274 61620 68280
rect 61580 63510 61608 68274
rect 61568 63504 61620 63510
rect 61568 63446 61620 63452
rect 64892 42158 64920 69414
rect 65064 69352 65116 69358
rect 65064 69294 65116 69300
rect 66352 69352 66404 69358
rect 66352 69294 66404 69300
rect 64972 69216 65024 69222
rect 64972 69158 65024 69164
rect 64984 68338 65012 69158
rect 64972 68332 65024 68338
rect 64972 68274 65024 68280
rect 65076 68270 65104 69294
rect 66260 69216 66312 69222
rect 66260 69158 66312 69164
rect 65654 69116 65962 69136
rect 65654 69114 65660 69116
rect 65716 69114 65740 69116
rect 65796 69114 65820 69116
rect 65876 69114 65900 69116
rect 65956 69114 65962 69116
rect 65716 69062 65718 69114
rect 65898 69062 65900 69114
rect 65654 69060 65660 69062
rect 65716 69060 65740 69062
rect 65796 69060 65820 69062
rect 65876 69060 65900 69062
rect 65956 69060 65962 69062
rect 65654 69040 65962 69060
rect 66272 68882 66300 69158
rect 66260 68876 66312 68882
rect 66260 68818 66312 68824
rect 65708 68672 65760 68678
rect 65708 68614 65760 68620
rect 65720 68406 65748 68614
rect 65708 68400 65760 68406
rect 65708 68342 65760 68348
rect 65064 68264 65116 68270
rect 65064 68206 65116 68212
rect 65654 68028 65962 68048
rect 65654 68026 65660 68028
rect 65716 68026 65740 68028
rect 65796 68026 65820 68028
rect 65876 68026 65900 68028
rect 65956 68026 65962 68028
rect 65716 67974 65718 68026
rect 65898 67974 65900 68026
rect 65654 67972 65660 67974
rect 65716 67972 65740 67974
rect 65796 67972 65820 67974
rect 65876 67972 65900 67974
rect 65956 67972 65962 67974
rect 65654 67952 65962 67972
rect 66364 67930 66392 69294
rect 67008 68270 67036 71200
rect 67730 70136 67786 70145
rect 67730 70071 67786 70080
rect 67088 68740 67140 68746
rect 67088 68682 67140 68688
rect 66996 68264 67048 68270
rect 66996 68206 67048 68212
rect 67100 67930 67128 68682
rect 67272 68196 67324 68202
rect 67272 68138 67324 68144
rect 66352 67924 66404 67930
rect 66352 67866 66404 67872
rect 67088 67924 67140 67930
rect 67088 67866 67140 67872
rect 66720 67720 66772 67726
rect 66720 67662 66772 67668
rect 65654 66940 65962 66960
rect 65654 66938 65660 66940
rect 65716 66938 65740 66940
rect 65796 66938 65820 66940
rect 65876 66938 65900 66940
rect 65956 66938 65962 66940
rect 65716 66886 65718 66938
rect 65898 66886 65900 66938
rect 65654 66884 65660 66886
rect 65716 66884 65740 66886
rect 65796 66884 65820 66886
rect 65876 66884 65900 66886
rect 65956 66884 65962 66886
rect 65654 66864 65962 66884
rect 65654 65852 65962 65872
rect 65654 65850 65660 65852
rect 65716 65850 65740 65852
rect 65796 65850 65820 65852
rect 65876 65850 65900 65852
rect 65956 65850 65962 65852
rect 65716 65798 65718 65850
rect 65898 65798 65900 65850
rect 65654 65796 65660 65798
rect 65716 65796 65740 65798
rect 65796 65796 65820 65798
rect 65876 65796 65900 65798
rect 65956 65796 65962 65798
rect 65654 65776 65962 65796
rect 65654 64764 65962 64784
rect 65654 64762 65660 64764
rect 65716 64762 65740 64764
rect 65796 64762 65820 64764
rect 65876 64762 65900 64764
rect 65956 64762 65962 64764
rect 65716 64710 65718 64762
rect 65898 64710 65900 64762
rect 65654 64708 65660 64710
rect 65716 64708 65740 64710
rect 65796 64708 65820 64710
rect 65876 64708 65900 64710
rect 65956 64708 65962 64710
rect 65654 64688 65962 64708
rect 66260 63776 66312 63782
rect 66260 63718 66312 63724
rect 65654 63676 65962 63696
rect 65654 63674 65660 63676
rect 65716 63674 65740 63676
rect 65796 63674 65820 63676
rect 65876 63674 65900 63676
rect 65956 63674 65962 63676
rect 65716 63622 65718 63674
rect 65898 63622 65900 63674
rect 65654 63620 65660 63622
rect 65716 63620 65740 63622
rect 65796 63620 65820 63622
rect 65876 63620 65900 63622
rect 65956 63620 65962 63622
rect 65654 63600 65962 63620
rect 66272 63442 66300 63718
rect 66260 63436 66312 63442
rect 66260 63378 66312 63384
rect 66444 63300 66496 63306
rect 66444 63242 66496 63248
rect 66456 63034 66484 63242
rect 66444 63028 66496 63034
rect 66444 62970 66496 62976
rect 65654 62588 65962 62608
rect 65654 62586 65660 62588
rect 65716 62586 65740 62588
rect 65796 62586 65820 62588
rect 65876 62586 65900 62588
rect 65956 62586 65962 62588
rect 65716 62534 65718 62586
rect 65898 62534 65900 62586
rect 65654 62532 65660 62534
rect 65716 62532 65740 62534
rect 65796 62532 65820 62534
rect 65876 62532 65900 62534
rect 65956 62532 65962 62534
rect 65654 62512 65962 62532
rect 66260 62280 66312 62286
rect 66260 62222 66312 62228
rect 66272 61878 66300 62222
rect 66260 61872 66312 61878
rect 66260 61814 66312 61820
rect 65654 61500 65962 61520
rect 65654 61498 65660 61500
rect 65716 61498 65740 61500
rect 65796 61498 65820 61500
rect 65876 61498 65900 61500
rect 65956 61498 65962 61500
rect 65716 61446 65718 61498
rect 65898 61446 65900 61498
rect 65654 61444 65660 61446
rect 65716 61444 65740 61446
rect 65796 61444 65820 61446
rect 65876 61444 65900 61446
rect 65956 61444 65962 61446
rect 65654 61424 65962 61444
rect 65654 60412 65962 60432
rect 65654 60410 65660 60412
rect 65716 60410 65740 60412
rect 65796 60410 65820 60412
rect 65876 60410 65900 60412
rect 65956 60410 65962 60412
rect 65716 60358 65718 60410
rect 65898 60358 65900 60410
rect 65654 60356 65660 60358
rect 65716 60356 65740 60358
rect 65796 60356 65820 60358
rect 65876 60356 65900 60358
rect 65956 60356 65962 60358
rect 65654 60336 65962 60356
rect 65654 59324 65962 59344
rect 65654 59322 65660 59324
rect 65716 59322 65740 59324
rect 65796 59322 65820 59324
rect 65876 59322 65900 59324
rect 65956 59322 65962 59324
rect 65716 59270 65718 59322
rect 65898 59270 65900 59322
rect 65654 59268 65660 59270
rect 65716 59268 65740 59270
rect 65796 59268 65820 59270
rect 65876 59268 65900 59270
rect 65956 59268 65962 59270
rect 65654 59248 65962 59268
rect 66260 58336 66312 58342
rect 66260 58278 66312 58284
rect 65654 58236 65962 58256
rect 65654 58234 65660 58236
rect 65716 58234 65740 58236
rect 65796 58234 65820 58236
rect 65876 58234 65900 58236
rect 65956 58234 65962 58236
rect 65716 58182 65718 58234
rect 65898 58182 65900 58234
rect 65654 58180 65660 58182
rect 65716 58180 65740 58182
rect 65796 58180 65820 58182
rect 65876 58180 65900 58182
rect 65956 58180 65962 58182
rect 65654 58160 65962 58180
rect 66272 57934 66300 58278
rect 66260 57928 66312 57934
rect 66260 57870 66312 57876
rect 66444 57860 66496 57866
rect 66444 57802 66496 57808
rect 66456 57594 66484 57802
rect 66444 57588 66496 57594
rect 66444 57530 66496 57536
rect 65654 57148 65962 57168
rect 65654 57146 65660 57148
rect 65716 57146 65740 57148
rect 65796 57146 65820 57148
rect 65876 57146 65900 57148
rect 65956 57146 65962 57148
rect 65716 57094 65718 57146
rect 65898 57094 65900 57146
rect 65654 57092 65660 57094
rect 65716 57092 65740 57094
rect 65796 57092 65820 57094
rect 65876 57092 65900 57094
rect 65956 57092 65962 57094
rect 65654 57072 65962 57092
rect 65654 56060 65962 56080
rect 65654 56058 65660 56060
rect 65716 56058 65740 56060
rect 65796 56058 65820 56060
rect 65876 56058 65900 56060
rect 65956 56058 65962 56060
rect 65716 56006 65718 56058
rect 65898 56006 65900 56058
rect 65654 56004 65660 56006
rect 65716 56004 65740 56006
rect 65796 56004 65820 56006
rect 65876 56004 65900 56006
rect 65956 56004 65962 56006
rect 65654 55984 65962 56004
rect 66166 55176 66222 55185
rect 66166 55111 66222 55120
rect 65654 54972 65962 54992
rect 65654 54970 65660 54972
rect 65716 54970 65740 54972
rect 65796 54970 65820 54972
rect 65876 54970 65900 54972
rect 65956 54970 65962 54972
rect 65716 54918 65718 54970
rect 65898 54918 65900 54970
rect 65654 54916 65660 54918
rect 65716 54916 65740 54918
rect 65796 54916 65820 54918
rect 65876 54916 65900 54918
rect 65956 54916 65962 54918
rect 65654 54896 65962 54916
rect 65654 53884 65962 53904
rect 65654 53882 65660 53884
rect 65716 53882 65740 53884
rect 65796 53882 65820 53884
rect 65876 53882 65900 53884
rect 65956 53882 65962 53884
rect 65716 53830 65718 53882
rect 65898 53830 65900 53882
rect 65654 53828 65660 53830
rect 65716 53828 65740 53830
rect 65796 53828 65820 53830
rect 65876 53828 65900 53830
rect 65956 53828 65962 53830
rect 65654 53808 65962 53828
rect 65654 52796 65962 52816
rect 65654 52794 65660 52796
rect 65716 52794 65740 52796
rect 65796 52794 65820 52796
rect 65876 52794 65900 52796
rect 65956 52794 65962 52796
rect 65716 52742 65718 52794
rect 65898 52742 65900 52794
rect 65654 52740 65660 52742
rect 65716 52740 65740 52742
rect 65796 52740 65820 52742
rect 65876 52740 65900 52742
rect 65956 52740 65962 52742
rect 65654 52720 65962 52740
rect 66076 51808 66128 51814
rect 66076 51750 66128 51756
rect 65654 51708 65962 51728
rect 65654 51706 65660 51708
rect 65716 51706 65740 51708
rect 65796 51706 65820 51708
rect 65876 51706 65900 51708
rect 65956 51706 65962 51708
rect 65716 51654 65718 51706
rect 65898 51654 65900 51706
rect 65654 51652 65660 51654
rect 65716 51652 65740 51654
rect 65796 51652 65820 51654
rect 65876 51652 65900 51654
rect 65956 51652 65962 51654
rect 65654 51632 65962 51652
rect 65654 50620 65962 50640
rect 65654 50618 65660 50620
rect 65716 50618 65740 50620
rect 65796 50618 65820 50620
rect 65876 50618 65900 50620
rect 65956 50618 65962 50620
rect 65716 50566 65718 50618
rect 65898 50566 65900 50618
rect 65654 50564 65660 50566
rect 65716 50564 65740 50566
rect 65796 50564 65820 50566
rect 65876 50564 65900 50566
rect 65956 50564 65962 50566
rect 65654 50544 65962 50564
rect 65522 49736 65578 49745
rect 65522 49671 65578 49680
rect 64880 42152 64932 42158
rect 64880 42094 64932 42100
rect 60740 41064 60792 41070
rect 60740 41006 60792 41012
rect 65536 32842 65564 49671
rect 65654 49532 65962 49552
rect 65654 49530 65660 49532
rect 65716 49530 65740 49532
rect 65796 49530 65820 49532
rect 65876 49530 65900 49532
rect 65956 49530 65962 49532
rect 65716 49478 65718 49530
rect 65898 49478 65900 49530
rect 65654 49476 65660 49478
rect 65716 49476 65740 49478
rect 65796 49476 65820 49478
rect 65876 49476 65900 49478
rect 65956 49476 65962 49478
rect 65654 49456 65962 49476
rect 65654 48444 65962 48464
rect 65654 48442 65660 48444
rect 65716 48442 65740 48444
rect 65796 48442 65820 48444
rect 65876 48442 65900 48444
rect 65956 48442 65962 48444
rect 65716 48390 65718 48442
rect 65898 48390 65900 48442
rect 65654 48388 65660 48390
rect 65716 48388 65740 48390
rect 65796 48388 65820 48390
rect 65876 48388 65900 48390
rect 65956 48388 65962 48390
rect 65654 48368 65962 48388
rect 65654 47356 65962 47376
rect 65654 47354 65660 47356
rect 65716 47354 65740 47356
rect 65796 47354 65820 47356
rect 65876 47354 65900 47356
rect 65956 47354 65962 47356
rect 65716 47302 65718 47354
rect 65898 47302 65900 47354
rect 65654 47300 65660 47302
rect 65716 47300 65740 47302
rect 65796 47300 65820 47302
rect 65876 47300 65900 47302
rect 65956 47300 65962 47302
rect 65654 47280 65962 47300
rect 65654 46268 65962 46288
rect 65654 46266 65660 46268
rect 65716 46266 65740 46268
rect 65796 46266 65820 46268
rect 65876 46266 65900 46268
rect 65956 46266 65962 46268
rect 65716 46214 65718 46266
rect 65898 46214 65900 46266
rect 65654 46212 65660 46214
rect 65716 46212 65740 46214
rect 65796 46212 65820 46214
rect 65876 46212 65900 46214
rect 65956 46212 65962 46214
rect 65654 46192 65962 46212
rect 65654 45180 65962 45200
rect 65654 45178 65660 45180
rect 65716 45178 65740 45180
rect 65796 45178 65820 45180
rect 65876 45178 65900 45180
rect 65956 45178 65962 45180
rect 65716 45126 65718 45178
rect 65898 45126 65900 45178
rect 65654 45124 65660 45126
rect 65716 45124 65740 45126
rect 65796 45124 65820 45126
rect 65876 45124 65900 45126
rect 65956 45124 65962 45126
rect 65654 45104 65962 45124
rect 65654 44092 65962 44112
rect 65654 44090 65660 44092
rect 65716 44090 65740 44092
rect 65796 44090 65820 44092
rect 65876 44090 65900 44092
rect 65956 44090 65962 44092
rect 65716 44038 65718 44090
rect 65898 44038 65900 44090
rect 65654 44036 65660 44038
rect 65716 44036 65740 44038
rect 65796 44036 65820 44038
rect 65876 44036 65900 44038
rect 65956 44036 65962 44038
rect 65654 44016 65962 44036
rect 65654 43004 65962 43024
rect 65654 43002 65660 43004
rect 65716 43002 65740 43004
rect 65796 43002 65820 43004
rect 65876 43002 65900 43004
rect 65956 43002 65962 43004
rect 65716 42950 65718 43002
rect 65898 42950 65900 43002
rect 65654 42948 65660 42950
rect 65716 42948 65740 42950
rect 65796 42948 65820 42950
rect 65876 42948 65900 42950
rect 65956 42948 65962 42950
rect 65654 42928 65962 42948
rect 65800 42696 65852 42702
rect 65800 42638 65852 42644
rect 65812 42226 65840 42638
rect 65800 42220 65852 42226
rect 65800 42162 65852 42168
rect 65984 42152 66036 42158
rect 65984 42094 66036 42100
rect 65654 41916 65962 41936
rect 65654 41914 65660 41916
rect 65716 41914 65740 41916
rect 65796 41914 65820 41916
rect 65876 41914 65900 41916
rect 65956 41914 65962 41916
rect 65716 41862 65718 41914
rect 65898 41862 65900 41914
rect 65654 41860 65660 41862
rect 65716 41860 65740 41862
rect 65796 41860 65820 41862
rect 65876 41860 65900 41862
rect 65956 41860 65962 41862
rect 65654 41840 65962 41860
rect 65996 41818 66024 42094
rect 65984 41812 66036 41818
rect 65984 41754 66036 41760
rect 66088 41698 66116 51750
rect 65996 41670 66116 41698
rect 65654 40828 65962 40848
rect 65654 40826 65660 40828
rect 65716 40826 65740 40828
rect 65796 40826 65820 40828
rect 65876 40826 65900 40828
rect 65956 40826 65962 40828
rect 65716 40774 65718 40826
rect 65898 40774 65900 40826
rect 65654 40772 65660 40774
rect 65716 40772 65740 40774
rect 65796 40772 65820 40774
rect 65876 40772 65900 40774
rect 65956 40772 65962 40774
rect 65654 40752 65962 40772
rect 65654 39740 65962 39760
rect 65654 39738 65660 39740
rect 65716 39738 65740 39740
rect 65796 39738 65820 39740
rect 65876 39738 65900 39740
rect 65956 39738 65962 39740
rect 65716 39686 65718 39738
rect 65898 39686 65900 39738
rect 65654 39684 65660 39686
rect 65716 39684 65740 39686
rect 65796 39684 65820 39686
rect 65876 39684 65900 39686
rect 65956 39684 65962 39686
rect 65654 39664 65962 39684
rect 65654 38652 65962 38672
rect 65654 38650 65660 38652
rect 65716 38650 65740 38652
rect 65796 38650 65820 38652
rect 65876 38650 65900 38652
rect 65956 38650 65962 38652
rect 65716 38598 65718 38650
rect 65898 38598 65900 38650
rect 65654 38596 65660 38598
rect 65716 38596 65740 38598
rect 65796 38596 65820 38598
rect 65876 38596 65900 38598
rect 65956 38596 65962 38598
rect 65654 38576 65962 38596
rect 65654 37564 65962 37584
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37488 65962 37508
rect 65654 36476 65962 36496
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36400 65962 36420
rect 65996 35894 66024 41670
rect 66180 41414 66208 55111
rect 66444 51332 66496 51338
rect 66444 51274 66496 51280
rect 66456 51066 66484 51274
rect 66444 51060 66496 51066
rect 66444 51002 66496 51008
rect 66260 47048 66312 47054
rect 66260 46990 66312 46996
rect 66272 46646 66300 46990
rect 66260 46640 66312 46646
rect 66260 46582 66312 46588
rect 66260 45280 66312 45286
rect 66260 45222 66312 45228
rect 66272 44946 66300 45222
rect 66260 44940 66312 44946
rect 66260 44882 66312 44888
rect 66444 44804 66496 44810
rect 66444 44746 66496 44752
rect 66456 44538 66484 44746
rect 66444 44532 66496 44538
rect 66444 44474 66496 44480
rect 66628 44396 66680 44402
rect 66628 44338 66680 44344
rect 66444 43716 66496 43722
rect 66444 43658 66496 43664
rect 66456 43450 66484 43658
rect 66444 43444 66496 43450
rect 66444 43386 66496 43392
rect 66088 41386 66208 41414
rect 66088 40118 66116 41386
rect 66260 40928 66312 40934
rect 66260 40870 66312 40876
rect 66272 40594 66300 40870
rect 66260 40588 66312 40594
rect 66260 40530 66312 40536
rect 66076 40112 66128 40118
rect 66076 40054 66128 40060
rect 66640 38214 66668 44338
rect 66628 38208 66680 38214
rect 66628 38150 66680 38156
rect 65996 35866 66116 35894
rect 65984 35624 66036 35630
rect 65984 35566 66036 35572
rect 65654 35388 65962 35408
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35312 65962 35332
rect 65996 35290 66024 35566
rect 65984 35284 66036 35290
rect 65984 35226 66036 35232
rect 65654 34300 65962 34320
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34224 65962 34244
rect 65654 33212 65962 33232
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33136 65962 33156
rect 65524 32836 65576 32842
rect 65524 32778 65576 32784
rect 65654 32124 65962 32144
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32048 65962 32068
rect 65984 31272 66036 31278
rect 65984 31214 66036 31220
rect 65654 31036 65962 31056
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30960 65962 30980
rect 65996 30938 66024 31214
rect 65984 30932 66036 30938
rect 65984 30874 66036 30880
rect 65654 29948 65962 29968
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29872 65962 29892
rect 65654 28860 65962 28880
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28784 65962 28804
rect 65654 27772 65962 27792
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27696 65962 27716
rect 65654 26684 65962 26704
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26608 65962 26628
rect 66088 26234 66116 35866
rect 66260 33312 66312 33318
rect 66260 33254 66312 33260
rect 66272 32978 66300 33254
rect 66260 32972 66312 32978
rect 66260 32914 66312 32920
rect 66444 32836 66496 32842
rect 66444 32778 66496 32784
rect 66456 32570 66484 32778
rect 66444 32564 66496 32570
rect 66444 32506 66496 32512
rect 66260 31816 66312 31822
rect 66260 31758 66312 31764
rect 66272 31414 66300 31758
rect 66260 31408 66312 31414
rect 66260 31350 66312 31356
rect 66168 30320 66220 30326
rect 66168 30262 66220 30268
rect 66180 30025 66208 30262
rect 66166 30016 66222 30025
rect 66166 29951 66222 29960
rect 65996 26206 66116 26234
rect 65654 25596 65962 25616
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25520 65962 25540
rect 65654 24508 65962 24528
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24432 65962 24452
rect 65654 23420 65962 23440
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23344 65962 23364
rect 65654 22332 65962 22352
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22256 65962 22276
rect 65996 21622 66024 26206
rect 66260 23520 66312 23526
rect 66260 23462 66312 23468
rect 66272 23186 66300 23462
rect 66260 23180 66312 23186
rect 66260 23122 66312 23128
rect 66444 23044 66496 23050
rect 66444 22986 66496 22992
rect 66456 22778 66484 22986
rect 66444 22772 66496 22778
rect 66444 22714 66496 22720
rect 66260 22160 66312 22166
rect 66260 22102 66312 22108
rect 65984 21616 66036 21622
rect 65984 21558 66036 21564
rect 66272 21486 66300 22102
rect 66260 21480 66312 21486
rect 66260 21422 66312 21428
rect 65654 21244 65962 21264
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21168 65962 21188
rect 65654 20156 65962 20176
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20080 65962 20100
rect 65654 19068 65962 19088
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 18992 65962 19012
rect 65654 17980 65962 18000
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17904 65962 17924
rect 65800 17672 65852 17678
rect 65800 17614 65852 17620
rect 65812 17202 65840 17614
rect 65800 17196 65852 17202
rect 65800 17138 65852 17144
rect 65654 16892 65962 16912
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16816 65962 16836
rect 66732 16658 66760 67662
rect 66996 67108 67048 67114
rect 66996 67050 67048 67056
rect 67008 66842 67036 67050
rect 66996 66836 67048 66842
rect 66996 66778 67048 66784
rect 66996 66020 67048 66026
rect 66996 65962 67048 65968
rect 67008 65754 67036 65962
rect 66996 65748 67048 65754
rect 66996 65690 67048 65696
rect 67284 65550 67312 68138
rect 67744 67726 67772 70071
rect 68296 69494 68324 71200
rect 68284 69488 68336 69494
rect 68284 69430 68336 69436
rect 69584 68882 69612 71200
rect 69572 68876 69624 68882
rect 69572 68818 69624 68824
rect 67732 67720 67784 67726
rect 67732 67662 67784 67668
rect 67638 67416 67694 67425
rect 67638 67351 67694 67360
rect 67652 67318 67680 67351
rect 67640 67312 67692 67318
rect 67640 67254 67692 67260
rect 67548 67176 67600 67182
rect 67548 67118 67600 67124
rect 67560 66842 67588 67118
rect 67548 66836 67600 66842
rect 67548 66778 67600 66784
rect 67456 66632 67508 66638
rect 67456 66574 67508 66580
rect 67364 66088 67416 66094
rect 67364 66030 67416 66036
rect 67376 65754 67404 66030
rect 67364 65748 67416 65754
rect 67364 65690 67416 65696
rect 67272 65544 67324 65550
rect 67272 65486 67324 65492
rect 67284 60058 67312 65486
rect 67364 60648 67416 60654
rect 67364 60590 67416 60596
rect 67376 60314 67404 60590
rect 67364 60308 67416 60314
rect 67364 60250 67416 60256
rect 67284 60030 67404 60058
rect 67272 59628 67324 59634
rect 67272 59570 67324 59576
rect 67180 59424 67232 59430
rect 67180 59366 67232 59372
rect 66996 57452 67048 57458
rect 66996 57394 67048 57400
rect 66812 50924 66864 50930
rect 66812 50866 66864 50872
rect 66824 46170 66852 50866
rect 67008 47122 67036 57394
rect 67088 56704 67140 56710
rect 67088 56646 67140 56652
rect 66996 47116 67048 47122
rect 66996 47058 67048 47064
rect 67100 46986 67128 56646
rect 67192 55214 67220 59366
rect 67284 59265 67312 59570
rect 67270 59256 67326 59265
rect 67270 59191 67326 59200
rect 67192 55186 67312 55214
rect 67180 47116 67232 47122
rect 67180 47058 67232 47064
rect 67088 46980 67140 46986
rect 67088 46922 67140 46928
rect 67192 46866 67220 47058
rect 67008 46838 67220 46866
rect 66812 46164 66864 46170
rect 66812 46106 66864 46112
rect 66812 45960 66864 45966
rect 66812 45902 66864 45908
rect 66824 38350 66852 45902
rect 67008 43314 67036 46838
rect 67284 46730 67312 55186
rect 67100 46702 67312 46730
rect 66996 43308 67048 43314
rect 66996 43250 67048 43256
rect 67008 41614 67036 43250
rect 67100 42362 67128 46702
rect 67376 46594 67404 60030
rect 67284 46566 67404 46594
rect 67180 46164 67232 46170
rect 67180 46106 67232 46112
rect 67088 42356 67140 42362
rect 67088 42298 67140 42304
rect 66996 41608 67048 41614
rect 66996 41550 67048 41556
rect 67088 40928 67140 40934
rect 67088 40870 67140 40876
rect 67100 40594 67128 40870
rect 67088 40588 67140 40594
rect 67088 40530 67140 40536
rect 66812 38344 66864 38350
rect 66812 38286 66864 38292
rect 66812 38208 66864 38214
rect 66812 38150 66864 38156
rect 66824 30734 66852 38150
rect 66904 36168 66956 36174
rect 66904 36110 66956 36116
rect 66916 35766 66944 36110
rect 66904 35760 66956 35766
rect 66904 35702 66956 35708
rect 66812 30728 66864 30734
rect 66812 30670 66864 30676
rect 67192 22642 67220 46106
rect 67284 41138 67312 46566
rect 67364 46504 67416 46510
rect 67364 46446 67416 46452
rect 67376 46170 67404 46446
rect 67364 46164 67416 46170
rect 67364 46106 67416 46112
rect 67272 41132 67324 41138
rect 67272 41074 67324 41080
rect 67272 40112 67324 40118
rect 67272 40054 67324 40060
rect 67284 39545 67312 40054
rect 67364 39840 67416 39846
rect 67364 39782 67416 39788
rect 67270 39536 67326 39545
rect 67270 39471 67326 39480
rect 67376 35834 67404 39782
rect 67364 35828 67416 35834
rect 67364 35770 67416 35776
rect 67468 35086 67496 66574
rect 67548 66088 67600 66094
rect 67546 66056 67548 66065
rect 67600 66056 67602 66065
rect 67546 65991 67602 66000
rect 68100 63368 68152 63374
rect 68098 63336 68100 63345
rect 68152 63336 68154 63345
rect 68098 63271 68154 63280
rect 67548 62892 67600 62898
rect 67548 62834 67600 62840
rect 67560 61198 67588 62834
rect 67638 61976 67694 61985
rect 67638 61911 67694 61920
rect 67652 61878 67680 61911
rect 67640 61872 67692 61878
rect 67640 61814 67692 61820
rect 67640 61736 67692 61742
rect 67640 61678 67692 61684
rect 67652 61402 67680 61678
rect 67640 61396 67692 61402
rect 67640 61338 67692 61344
rect 67548 61192 67600 61198
rect 67548 61134 67600 61140
rect 67548 60648 67600 60654
rect 67546 60616 67548 60625
rect 67600 60616 67602 60625
rect 67546 60551 67602 60560
rect 68100 60580 68152 60586
rect 68100 60522 68152 60528
rect 68112 60314 68140 60522
rect 68100 60308 68152 60314
rect 68100 60250 68152 60256
rect 68100 57928 68152 57934
rect 68098 57896 68100 57905
rect 68152 57896 68154 57905
rect 68098 57831 68154 57840
rect 67548 56840 67600 56846
rect 67548 56782 67600 56788
rect 67560 56545 67588 56782
rect 67546 56536 67602 56545
rect 67546 56471 67602 56480
rect 68100 51332 68152 51338
rect 68100 51274 68152 51280
rect 68112 51105 68140 51274
rect 68098 51096 68154 51105
rect 68098 51031 68154 51040
rect 67732 48068 67784 48074
rect 67732 48010 67784 48016
rect 67744 47705 67772 48010
rect 67824 48000 67876 48006
rect 67824 47942 67876 47948
rect 67836 47802 67864 47942
rect 67824 47796 67876 47802
rect 67824 47738 67876 47744
rect 67730 47696 67786 47705
rect 67730 47631 67786 47640
rect 67548 46504 67600 46510
rect 67548 46446 67600 46452
rect 67560 46345 67588 46446
rect 67546 46336 67602 46345
rect 67546 46271 67602 46280
rect 68098 44976 68154 44985
rect 68098 44911 68100 44920
rect 68152 44911 68154 44920
rect 68100 44882 68152 44888
rect 67916 43852 67968 43858
rect 67916 43794 67968 43800
rect 67928 42770 67956 43794
rect 68100 43716 68152 43722
rect 68100 43658 68152 43664
rect 68112 43625 68140 43658
rect 68098 43616 68154 43625
rect 68098 43551 68154 43560
rect 67916 42764 67968 42770
rect 67916 42706 67968 42712
rect 67546 42256 67602 42265
rect 67546 42191 67602 42200
rect 67560 42158 67588 42191
rect 67548 42152 67600 42158
rect 67548 42094 67600 42100
rect 68098 40896 68154 40905
rect 68098 40831 68154 40840
rect 68112 40594 68140 40831
rect 68100 40588 68152 40594
rect 68100 40530 68152 40536
rect 67548 35624 67600 35630
rect 67548 35566 67600 35572
rect 67560 35465 67588 35566
rect 67546 35456 67602 35465
rect 67546 35391 67602 35400
rect 67456 35080 67508 35086
rect 67456 35022 67508 35028
rect 67272 34604 67324 34610
rect 67272 34546 67324 34552
rect 67284 34105 67312 34546
rect 67270 34096 67326 34105
rect 67270 34031 67326 34040
rect 67272 33040 67324 33046
rect 67272 32982 67324 32988
rect 67284 32434 67312 32982
rect 67272 32428 67324 32434
rect 67272 32370 67324 32376
rect 67180 22636 67232 22642
rect 67180 22578 67232 22584
rect 66720 16652 66772 16658
rect 66720 16594 66772 16600
rect 66168 16584 66220 16590
rect 66168 16526 66220 16532
rect 65654 15804 65962 15824
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15728 65962 15748
rect 66180 15745 66208 16526
rect 66166 15736 66222 15745
rect 66166 15671 66222 15680
rect 66260 15360 66312 15366
rect 66260 15302 66312 15308
rect 66272 15094 66300 15302
rect 66260 15088 66312 15094
rect 66260 15030 66312 15036
rect 65654 14716 65962 14736
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14640 65962 14660
rect 65654 13628 65962 13648
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13552 65962 13572
rect 65654 12540 65962 12560
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12464 65962 12484
rect 65654 11452 65962 11472
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11376 65962 11396
rect 65654 10364 65962 10384
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10288 65962 10308
rect 65654 9276 65962 9296
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9200 65962 9220
rect 65654 8188 65962 8208
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8112 65962 8132
rect 65654 7100 65962 7120
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7024 65962 7044
rect 67192 6914 67220 22578
rect 67284 15502 67312 32370
rect 67272 15496 67324 15502
rect 67272 15438 67324 15444
rect 67364 14952 67416 14958
rect 67364 14894 67416 14900
rect 67376 14618 67404 14894
rect 67364 14612 67416 14618
rect 67364 14554 67416 14560
rect 67468 11778 67496 35022
rect 68100 32836 68152 32842
rect 68100 32778 68152 32784
rect 68112 32745 68140 32778
rect 68098 32736 68154 32745
rect 68098 32671 68154 32680
rect 67546 31376 67602 31385
rect 67546 31311 67602 31320
rect 67560 31278 67588 31311
rect 67548 31272 67600 31278
rect 67548 31214 67600 31220
rect 67548 30728 67600 30734
rect 67548 30670 67600 30676
rect 67560 21570 67588 30670
rect 68098 23216 68154 23225
rect 68098 23151 68100 23160
rect 68152 23151 68154 23160
rect 68100 23122 68152 23128
rect 67560 21542 67680 21570
rect 67548 21480 67600 21486
rect 67548 21422 67600 21428
rect 67560 21185 67588 21422
rect 67546 21176 67602 21185
rect 67546 21111 67602 21120
rect 67652 21026 67680 21542
rect 67560 20998 67680 21026
rect 67560 17218 67588 20998
rect 67824 18760 67876 18766
rect 67824 18702 67876 18708
rect 67836 18465 67864 18702
rect 68008 18624 68060 18630
rect 68008 18566 68060 18572
rect 67822 18456 67878 18465
rect 67822 18391 67878 18400
rect 68020 18290 68048 18566
rect 68008 18284 68060 18290
rect 68008 18226 68060 18232
rect 67732 17264 67784 17270
rect 67560 17190 67680 17218
rect 67732 17206 67784 17212
rect 67548 17128 67600 17134
rect 67546 17096 67548 17105
rect 67600 17096 67602 17105
rect 67546 17031 67602 17040
rect 67652 16946 67680 17190
rect 67560 16918 67680 16946
rect 67560 15042 67588 16918
rect 67744 16454 67772 17206
rect 67732 16448 67784 16454
rect 67732 16390 67784 16396
rect 67560 15014 67680 15042
rect 67548 14952 67600 14958
rect 67548 14894 67600 14900
rect 67560 14385 67588 14894
rect 67546 14376 67602 14385
rect 67546 14311 67602 14320
rect 67652 14226 67680 15014
rect 67100 6886 67220 6914
rect 67284 11750 67496 11778
rect 67560 14198 67680 14226
rect 65800 6792 65852 6798
rect 65800 6734 65852 6740
rect 65812 6322 65840 6734
rect 65800 6316 65852 6322
rect 65800 6258 65852 6264
rect 65984 6248 66036 6254
rect 65984 6190 66036 6196
rect 65654 6012 65962 6032
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5936 65962 5956
rect 65996 5914 66024 6190
rect 65984 5908 66036 5914
rect 65984 5850 66036 5856
rect 66444 5704 66496 5710
rect 66444 5646 66496 5652
rect 66456 5166 66484 5646
rect 66996 5568 67048 5574
rect 66996 5510 67048 5516
rect 67008 5302 67036 5510
rect 66996 5296 67048 5302
rect 66996 5238 67048 5244
rect 66444 5160 66496 5166
rect 66444 5102 66496 5108
rect 65654 4924 65962 4944
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4848 65962 4868
rect 66904 4616 66956 4622
rect 66904 4558 66956 4564
rect 66916 4010 66944 4558
rect 66904 4004 66956 4010
rect 66904 3946 66956 3952
rect 60648 3936 60700 3942
rect 60648 3878 60700 3884
rect 62120 3936 62172 3942
rect 62120 3878 62172 3884
rect 50896 3528 50948 3534
rect 50896 3470 50948 3476
rect 51724 3528 51776 3534
rect 51724 3470 51776 3476
rect 59728 3528 59780 3534
rect 59728 3470 59780 3476
rect 50620 1352 50672 1358
rect 50620 1294 50672 1300
rect 50908 800 50936 3470
rect 60660 3058 60688 3878
rect 62132 3602 62160 3878
rect 65654 3836 65962 3856
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3760 65962 3780
rect 62120 3596 62172 3602
rect 62120 3538 62172 3544
rect 62488 3596 62540 3602
rect 62488 3538 62540 3544
rect 62120 3460 62172 3466
rect 62120 3402 62172 3408
rect 60832 3392 60884 3398
rect 60832 3334 60884 3340
rect 60844 3126 60872 3334
rect 60832 3120 60884 3126
rect 60832 3062 60884 3068
rect 60648 3052 60700 3058
rect 60648 2994 60700 3000
rect 61200 2984 61252 2990
rect 61200 2926 61252 2932
rect 56048 2440 56100 2446
rect 56048 2382 56100 2388
rect 56060 800 56088 2382
rect 56416 2372 56468 2378
rect 56416 2314 56468 2320
rect 56428 2038 56456 2314
rect 56416 2032 56468 2038
rect 56416 1974 56468 1980
rect 61212 800 61240 2926
rect 62132 2650 62160 3402
rect 62120 2644 62172 2650
rect 62120 2586 62172 2592
rect 62500 800 62528 3538
rect 65800 3528 65852 3534
rect 65800 3470 65852 3476
rect 65812 3058 65840 3470
rect 65984 3392 66036 3398
rect 65984 3334 66036 3340
rect 65996 3126 66024 3334
rect 65984 3120 66036 3126
rect 65984 3062 66036 3068
rect 65800 3052 65852 3058
rect 65800 2994 65852 3000
rect 67100 2922 67128 6886
rect 67284 5794 67312 11750
rect 67560 6914 67588 14198
rect 67824 13320 67876 13326
rect 67824 13262 67876 13268
rect 67836 13025 67864 13262
rect 68008 13184 68060 13190
rect 68008 13126 68060 13132
rect 67822 13016 67878 13025
rect 67822 12951 67878 12960
rect 68020 12782 68048 13126
rect 68008 12776 68060 12782
rect 68008 12718 68060 12724
rect 67640 7880 67692 7886
rect 67640 7822 67692 7828
rect 67652 7585 67680 7822
rect 67638 7576 67694 7585
rect 67638 7511 67694 7520
rect 67192 5766 67312 5794
rect 67376 6886 67588 6914
rect 67192 3942 67220 5766
rect 67272 5704 67324 5710
rect 67272 5646 67324 5652
rect 67284 4622 67312 5646
rect 67272 4616 67324 4622
rect 67272 4558 67324 4564
rect 67180 3936 67232 3942
rect 67180 3878 67232 3884
rect 67376 3534 67404 6886
rect 67548 6248 67600 6254
rect 67546 6216 67548 6225
rect 67600 6216 67602 6225
rect 67546 6151 67602 6160
rect 67548 5160 67600 5166
rect 67548 5102 67600 5108
rect 67560 4865 67588 5102
rect 67546 4856 67602 4865
rect 67546 4791 67602 4800
rect 67456 4480 67508 4486
rect 67456 4422 67508 4428
rect 67468 4078 67496 4422
rect 67456 4072 67508 4078
rect 67456 4014 67508 4020
rect 68928 4072 68980 4078
rect 68928 4014 68980 4020
rect 67364 3528 67416 3534
rect 67364 3470 67416 3476
rect 67088 2916 67140 2922
rect 67088 2858 67140 2864
rect 65654 2748 65962 2768
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2672 65962 2692
rect 65064 2440 65116 2446
rect 65064 2382 65116 2388
rect 65076 800 65104 2382
rect 67640 2372 67692 2378
rect 67640 2314 67692 2320
rect 66168 1352 66220 1358
rect 66168 1294 66220 1300
rect 39500 734 39804 762
rect 39918 0 40030 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43782 0 43894 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 47002 0 47114 800
rect 48290 0 48402 800
rect 49578 0 49690 800
rect 50866 0 50978 800
rect 52154 0 52266 800
rect 53442 0 53554 800
rect 54730 0 54842 800
rect 56018 0 56130 800
rect 57306 0 57418 800
rect 58594 0 58706 800
rect 59882 0 59994 800
rect 61170 0 61282 800
rect 62458 0 62570 800
rect 63746 0 63858 800
rect 65034 0 65146 800
rect 66180 785 66208 1294
rect 67652 800 67680 2314
rect 68940 800 68968 4014
rect 69572 2984 69624 2990
rect 69572 2926 69624 2932
rect 69584 800 69612 2926
rect 66166 776 66222 785
rect 66166 711 66222 720
rect 66322 0 66434 800
rect 67610 0 67722 800
rect 68898 0 69010 800
rect 69542 0 69654 800
<< via2 >>
rect 1398 70896 1454 70952
rect 2778 68720 2834 68776
rect 1398 63316 1400 63336
rect 1400 63316 1452 63336
rect 1452 63316 1454 63336
rect 1398 63280 1454 63316
rect 1858 60560 1914 60616
rect 1398 56480 1454 56536
rect 1858 52400 1914 52456
rect 2778 67360 2834 67416
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 2778 59200 2834 59256
rect 2778 53760 2834 53816
rect 2778 47640 2834 47696
rect 1858 46280 1914 46336
rect 1858 44920 1914 44976
rect 1858 43560 1914 43616
rect 1858 42200 1914 42256
rect 2042 42200 2098 42256
rect 2778 39500 2834 39536
rect 2778 39480 2780 39500
rect 2780 39480 2832 39500
rect 2832 39480 2834 39500
rect 3238 40840 3294 40896
rect 3238 38120 3294 38176
rect 3238 36760 3294 36816
rect 2778 35400 2834 35456
rect 1398 34040 1454 34096
rect 2778 31320 2834 31376
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 1858 24520 1914 24576
rect 1858 21120 1914 21176
rect 1858 7520 1914 7576
rect 2870 29960 2926 30016
rect 3054 27240 3110 27296
rect 2778 25880 2834 25936
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 3514 55120 3570 55176
rect 3514 51040 3570 51096
rect 3514 49680 3570 49736
rect 2778 23840 2834 23896
rect 2778 22516 2780 22536
rect 2780 22516 2832 22536
rect 2832 22516 2834 22536
rect 2778 22480 2834 22516
rect 2962 15680 3018 15736
rect 2778 12960 2834 13016
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 3606 4800 3662 4856
rect 3146 3440 3202 3496
rect 2778 2080 2834 2136
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 19580 69658 19636 69660
rect 19660 69658 19716 69660
rect 19740 69658 19796 69660
rect 19820 69658 19876 69660
rect 19580 69606 19626 69658
rect 19626 69606 19636 69658
rect 19660 69606 19690 69658
rect 19690 69606 19702 69658
rect 19702 69606 19716 69658
rect 19740 69606 19754 69658
rect 19754 69606 19766 69658
rect 19766 69606 19796 69658
rect 19820 69606 19830 69658
rect 19830 69606 19876 69658
rect 19580 69604 19636 69606
rect 19660 69604 19716 69606
rect 19740 69604 19796 69606
rect 19820 69604 19876 69606
rect 19580 68570 19636 68572
rect 19660 68570 19716 68572
rect 19740 68570 19796 68572
rect 19820 68570 19876 68572
rect 19580 68518 19626 68570
rect 19626 68518 19636 68570
rect 19660 68518 19690 68570
rect 19690 68518 19702 68570
rect 19702 68518 19716 68570
rect 19740 68518 19754 68570
rect 19754 68518 19766 68570
rect 19766 68518 19796 68570
rect 19820 68518 19830 68570
rect 19830 68518 19876 68570
rect 19580 68516 19636 68518
rect 19660 68516 19716 68518
rect 19740 68516 19796 68518
rect 19820 68516 19876 68518
rect 19580 67482 19636 67484
rect 19660 67482 19716 67484
rect 19740 67482 19796 67484
rect 19820 67482 19876 67484
rect 19580 67430 19626 67482
rect 19626 67430 19636 67482
rect 19660 67430 19690 67482
rect 19690 67430 19702 67482
rect 19702 67430 19716 67482
rect 19740 67430 19754 67482
rect 19754 67430 19766 67482
rect 19766 67430 19796 67482
rect 19820 67430 19830 67482
rect 19830 67430 19876 67482
rect 19580 67428 19636 67430
rect 19660 67428 19716 67430
rect 19740 67428 19796 67430
rect 19820 67428 19876 67430
rect 19580 66394 19636 66396
rect 19660 66394 19716 66396
rect 19740 66394 19796 66396
rect 19820 66394 19876 66396
rect 19580 66342 19626 66394
rect 19626 66342 19636 66394
rect 19660 66342 19690 66394
rect 19690 66342 19702 66394
rect 19702 66342 19716 66394
rect 19740 66342 19754 66394
rect 19754 66342 19766 66394
rect 19766 66342 19796 66394
rect 19820 66342 19830 66394
rect 19830 66342 19876 66394
rect 19580 66340 19636 66342
rect 19660 66340 19716 66342
rect 19740 66340 19796 66342
rect 19820 66340 19876 66342
rect 19580 65306 19636 65308
rect 19660 65306 19716 65308
rect 19740 65306 19796 65308
rect 19820 65306 19876 65308
rect 19580 65254 19626 65306
rect 19626 65254 19636 65306
rect 19660 65254 19690 65306
rect 19690 65254 19702 65306
rect 19702 65254 19716 65306
rect 19740 65254 19754 65306
rect 19754 65254 19766 65306
rect 19766 65254 19796 65306
rect 19820 65254 19830 65306
rect 19830 65254 19876 65306
rect 19580 65252 19636 65254
rect 19660 65252 19716 65254
rect 19740 65252 19796 65254
rect 19820 65252 19876 65254
rect 19580 64218 19636 64220
rect 19660 64218 19716 64220
rect 19740 64218 19796 64220
rect 19820 64218 19876 64220
rect 19580 64166 19626 64218
rect 19626 64166 19636 64218
rect 19660 64166 19690 64218
rect 19690 64166 19702 64218
rect 19702 64166 19716 64218
rect 19740 64166 19754 64218
rect 19754 64166 19766 64218
rect 19766 64166 19796 64218
rect 19820 64166 19830 64218
rect 19830 64166 19876 64218
rect 19580 64164 19636 64166
rect 19660 64164 19716 64166
rect 19740 64164 19796 64166
rect 19820 64164 19876 64166
rect 19580 63130 19636 63132
rect 19660 63130 19716 63132
rect 19740 63130 19796 63132
rect 19820 63130 19876 63132
rect 19580 63078 19626 63130
rect 19626 63078 19636 63130
rect 19660 63078 19690 63130
rect 19690 63078 19702 63130
rect 19702 63078 19716 63130
rect 19740 63078 19754 63130
rect 19754 63078 19766 63130
rect 19766 63078 19796 63130
rect 19820 63078 19830 63130
rect 19830 63078 19876 63130
rect 19580 63076 19636 63078
rect 19660 63076 19716 63078
rect 19740 63076 19796 63078
rect 19820 63076 19876 63078
rect 19580 62042 19636 62044
rect 19660 62042 19716 62044
rect 19740 62042 19796 62044
rect 19820 62042 19876 62044
rect 19580 61990 19626 62042
rect 19626 61990 19636 62042
rect 19660 61990 19690 62042
rect 19690 61990 19702 62042
rect 19702 61990 19716 62042
rect 19740 61990 19754 62042
rect 19754 61990 19766 62042
rect 19766 61990 19796 62042
rect 19820 61990 19830 62042
rect 19830 61990 19876 62042
rect 19580 61988 19636 61990
rect 19660 61988 19716 61990
rect 19740 61988 19796 61990
rect 19820 61988 19876 61990
rect 19580 60954 19636 60956
rect 19660 60954 19716 60956
rect 19740 60954 19796 60956
rect 19820 60954 19876 60956
rect 19580 60902 19626 60954
rect 19626 60902 19636 60954
rect 19660 60902 19690 60954
rect 19690 60902 19702 60954
rect 19702 60902 19716 60954
rect 19740 60902 19754 60954
rect 19754 60902 19766 60954
rect 19766 60902 19796 60954
rect 19820 60902 19830 60954
rect 19830 60902 19876 60954
rect 19580 60900 19636 60902
rect 19660 60900 19716 60902
rect 19740 60900 19796 60902
rect 19820 60900 19876 60902
rect 19580 59866 19636 59868
rect 19660 59866 19716 59868
rect 19740 59866 19796 59868
rect 19820 59866 19876 59868
rect 19580 59814 19626 59866
rect 19626 59814 19636 59866
rect 19660 59814 19690 59866
rect 19690 59814 19702 59866
rect 19702 59814 19716 59866
rect 19740 59814 19754 59866
rect 19754 59814 19766 59866
rect 19766 59814 19796 59866
rect 19820 59814 19830 59866
rect 19830 59814 19876 59866
rect 19580 59812 19636 59814
rect 19660 59812 19716 59814
rect 19740 59812 19796 59814
rect 19820 59812 19876 59814
rect 19580 58778 19636 58780
rect 19660 58778 19716 58780
rect 19740 58778 19796 58780
rect 19820 58778 19876 58780
rect 19580 58726 19626 58778
rect 19626 58726 19636 58778
rect 19660 58726 19690 58778
rect 19690 58726 19702 58778
rect 19702 58726 19716 58778
rect 19740 58726 19754 58778
rect 19754 58726 19766 58778
rect 19766 58726 19796 58778
rect 19820 58726 19830 58778
rect 19830 58726 19876 58778
rect 19580 58724 19636 58726
rect 19660 58724 19716 58726
rect 19740 58724 19796 58726
rect 19820 58724 19876 58726
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4618 3440 4674 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 13542 3576 13598 3632
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 21178 41556 21180 41576
rect 21180 41556 21232 41576
rect 21232 41556 21234 41576
rect 21178 41520 21234 41556
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 22466 41520 22522 41576
rect 25870 49680 25926 49736
rect 26146 57996 26202 58032
rect 26146 57976 26148 57996
rect 26148 57976 26200 57996
rect 26200 57976 26202 57996
rect 34940 69114 34996 69116
rect 35020 69114 35076 69116
rect 35100 69114 35156 69116
rect 35180 69114 35236 69116
rect 34940 69062 34986 69114
rect 34986 69062 34996 69114
rect 35020 69062 35050 69114
rect 35050 69062 35062 69114
rect 35062 69062 35076 69114
rect 35100 69062 35114 69114
rect 35114 69062 35126 69114
rect 35126 69062 35156 69114
rect 35180 69062 35190 69114
rect 35190 69062 35236 69114
rect 34940 69060 34996 69062
rect 35020 69060 35076 69062
rect 35100 69060 35156 69062
rect 35180 69060 35236 69062
rect 34940 68026 34996 68028
rect 35020 68026 35076 68028
rect 35100 68026 35156 68028
rect 35180 68026 35236 68028
rect 34940 67974 34986 68026
rect 34986 67974 34996 68026
rect 35020 67974 35050 68026
rect 35050 67974 35062 68026
rect 35062 67974 35076 68026
rect 35100 67974 35114 68026
rect 35114 67974 35126 68026
rect 35126 67974 35156 68026
rect 35180 67974 35190 68026
rect 35190 67974 35236 68026
rect 34940 67972 34996 67974
rect 35020 67972 35076 67974
rect 35100 67972 35156 67974
rect 35180 67972 35236 67974
rect 34940 66938 34996 66940
rect 35020 66938 35076 66940
rect 35100 66938 35156 66940
rect 35180 66938 35236 66940
rect 34940 66886 34986 66938
rect 34986 66886 34996 66938
rect 35020 66886 35050 66938
rect 35050 66886 35062 66938
rect 35062 66886 35076 66938
rect 35100 66886 35114 66938
rect 35114 66886 35126 66938
rect 35126 66886 35156 66938
rect 35180 66886 35190 66938
rect 35190 66886 35236 66938
rect 34940 66884 34996 66886
rect 35020 66884 35076 66886
rect 35100 66884 35156 66886
rect 35180 66884 35236 66886
rect 34940 65850 34996 65852
rect 35020 65850 35076 65852
rect 35100 65850 35156 65852
rect 35180 65850 35236 65852
rect 34940 65798 34986 65850
rect 34986 65798 34996 65850
rect 35020 65798 35050 65850
rect 35050 65798 35062 65850
rect 35062 65798 35076 65850
rect 35100 65798 35114 65850
rect 35114 65798 35126 65850
rect 35126 65798 35156 65850
rect 35180 65798 35190 65850
rect 35190 65798 35236 65850
rect 34940 65796 34996 65798
rect 35020 65796 35076 65798
rect 35100 65796 35156 65798
rect 35180 65796 35236 65798
rect 34940 64762 34996 64764
rect 35020 64762 35076 64764
rect 35100 64762 35156 64764
rect 35180 64762 35236 64764
rect 34940 64710 34986 64762
rect 34986 64710 34996 64762
rect 35020 64710 35050 64762
rect 35050 64710 35062 64762
rect 35062 64710 35076 64762
rect 35100 64710 35114 64762
rect 35114 64710 35126 64762
rect 35126 64710 35156 64762
rect 35180 64710 35190 64762
rect 35190 64710 35236 64762
rect 34940 64708 34996 64710
rect 35020 64708 35076 64710
rect 35100 64708 35156 64710
rect 35180 64708 35236 64710
rect 26054 46452 26056 46472
rect 26056 46452 26108 46472
rect 26108 46452 26110 46472
rect 26054 46416 26110 46452
rect 26146 42220 26202 42256
rect 26146 42200 26148 42220
rect 26148 42200 26200 42220
rect 26200 42200 26202 42220
rect 26330 46436 26386 46472
rect 26330 46416 26332 46436
rect 26332 46416 26384 46436
rect 26384 46416 26386 46436
rect 28170 41556 28172 41576
rect 28172 41556 28224 41576
rect 28224 41556 28226 41576
rect 28170 41520 28226 41556
rect 30286 48048 30342 48104
rect 34940 63674 34996 63676
rect 35020 63674 35076 63676
rect 35100 63674 35156 63676
rect 35180 63674 35236 63676
rect 34940 63622 34986 63674
rect 34986 63622 34996 63674
rect 35020 63622 35050 63674
rect 35050 63622 35062 63674
rect 35062 63622 35076 63674
rect 35100 63622 35114 63674
rect 35114 63622 35126 63674
rect 35126 63622 35156 63674
rect 35180 63622 35190 63674
rect 35190 63622 35236 63674
rect 34940 63620 34996 63622
rect 35020 63620 35076 63622
rect 35100 63620 35156 63622
rect 35180 63620 35236 63622
rect 34940 62586 34996 62588
rect 35020 62586 35076 62588
rect 35100 62586 35156 62588
rect 35180 62586 35236 62588
rect 34940 62534 34986 62586
rect 34986 62534 34996 62586
rect 35020 62534 35050 62586
rect 35050 62534 35062 62586
rect 35062 62534 35076 62586
rect 35100 62534 35114 62586
rect 35114 62534 35126 62586
rect 35126 62534 35156 62586
rect 35180 62534 35190 62586
rect 35190 62534 35236 62586
rect 34940 62532 34996 62534
rect 35020 62532 35076 62534
rect 35100 62532 35156 62534
rect 35180 62532 35236 62534
rect 34940 61498 34996 61500
rect 35020 61498 35076 61500
rect 35100 61498 35156 61500
rect 35180 61498 35236 61500
rect 34940 61446 34986 61498
rect 34986 61446 34996 61498
rect 35020 61446 35050 61498
rect 35050 61446 35062 61498
rect 35062 61446 35076 61498
rect 35100 61446 35114 61498
rect 35114 61446 35126 61498
rect 35126 61446 35156 61498
rect 35180 61446 35190 61498
rect 35190 61446 35236 61498
rect 34940 61444 34996 61446
rect 35020 61444 35076 61446
rect 35100 61444 35156 61446
rect 35180 61444 35236 61446
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 34940 59322 34996 59324
rect 35020 59322 35076 59324
rect 35100 59322 35156 59324
rect 35180 59322 35236 59324
rect 34940 59270 34986 59322
rect 34986 59270 34996 59322
rect 35020 59270 35050 59322
rect 35050 59270 35062 59322
rect 35062 59270 35076 59322
rect 35100 59270 35114 59322
rect 35114 59270 35126 59322
rect 35126 59270 35156 59322
rect 35180 59270 35190 59322
rect 35190 59270 35236 59322
rect 34940 59268 34996 59270
rect 35020 59268 35076 59270
rect 35100 59268 35156 59270
rect 35180 59268 35236 59270
rect 34940 58234 34996 58236
rect 35020 58234 35076 58236
rect 35100 58234 35156 58236
rect 35180 58234 35236 58236
rect 34940 58182 34986 58234
rect 34986 58182 34996 58234
rect 35020 58182 35050 58234
rect 35050 58182 35062 58234
rect 35062 58182 35076 58234
rect 35100 58182 35114 58234
rect 35114 58182 35126 58234
rect 35126 58182 35156 58234
rect 35180 58182 35190 58234
rect 35190 58182 35236 58234
rect 34940 58180 34996 58182
rect 35020 58180 35076 58182
rect 35100 58180 35156 58182
rect 35180 58180 35236 58182
rect 32954 48220 32956 48240
rect 32956 48220 33008 48240
rect 33008 48220 33010 48240
rect 32954 48184 33010 48220
rect 33230 47912 33286 47968
rect 33966 48204 34022 48240
rect 33966 48184 33968 48204
rect 33968 48184 34020 48204
rect 34020 48184 34022 48204
rect 33874 47912 33930 47968
rect 33782 47796 33838 47832
rect 33782 47776 33784 47796
rect 33784 47776 33836 47796
rect 33836 47776 33838 47796
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34610 49272 34666 49328
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34886 49272 34942 49328
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 35990 47796 36046 47832
rect 35990 47776 35992 47796
rect 35992 47776 36044 47796
rect 36044 47776 36046 47796
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 32310 36624 32366 36680
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34886 36660 34888 36680
rect 34888 36660 34940 36680
rect 34940 36660 34942 36680
rect 34886 36624 34942 36660
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 36358 48048 36414 48104
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35622 35128 35678 35184
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35622 34720 35678 34776
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 37278 41692 37280 41712
rect 37280 41692 37332 41712
rect 37332 41692 37334 41712
rect 37278 41656 37334 41692
rect 37646 41792 37702 41848
rect 37646 41384 37702 41440
rect 38106 41540 38162 41576
rect 38106 41520 38108 41540
rect 38108 41520 38160 41540
rect 38160 41520 38162 41540
rect 38658 41112 38714 41168
rect 39026 41692 39028 41712
rect 39028 41692 39080 41712
rect 39080 41692 39082 41712
rect 39026 41656 39082 41692
rect 41418 52980 41420 53000
rect 41420 52980 41472 53000
rect 41472 52980 41474 53000
rect 41418 52944 41474 52980
rect 42706 52944 42762 53000
rect 42614 50904 42670 50960
rect 43902 50924 43958 50960
rect 43902 50904 43904 50924
rect 43904 50904 43956 50924
rect 43956 50904 43958 50924
rect 43718 49136 43774 49192
rect 38750 37884 38752 37904
rect 38752 37884 38804 37904
rect 38804 37884 38806 37904
rect 38750 37848 38806 37884
rect 39946 37884 39948 37904
rect 39948 37884 40000 37904
rect 40000 37884 40002 37904
rect 39946 37848 40002 37884
rect 40314 40976 40370 41032
rect 45650 49172 45652 49192
rect 45652 49172 45704 49192
rect 45704 49172 45706 49192
rect 45650 49136 45706 49172
rect 42246 41792 42302 41848
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 46386 40996 46442 41032
rect 46386 40976 46388 40996
rect 46388 40976 46440 40996
rect 46440 40976 46442 40996
rect 45650 39380 45652 39400
rect 45652 39380 45704 39400
rect 45704 39380 45706 39400
rect 45650 39344 45706 39380
rect 46754 39344 46810 39400
rect 50300 69658 50356 69660
rect 50380 69658 50436 69660
rect 50460 69658 50516 69660
rect 50540 69658 50596 69660
rect 50300 69606 50346 69658
rect 50346 69606 50356 69658
rect 50380 69606 50410 69658
rect 50410 69606 50422 69658
rect 50422 69606 50436 69658
rect 50460 69606 50474 69658
rect 50474 69606 50486 69658
rect 50486 69606 50516 69658
rect 50540 69606 50550 69658
rect 50550 69606 50596 69658
rect 50300 69604 50356 69606
rect 50380 69604 50436 69606
rect 50460 69604 50516 69606
rect 50540 69604 50596 69606
rect 50300 68570 50356 68572
rect 50380 68570 50436 68572
rect 50460 68570 50516 68572
rect 50540 68570 50596 68572
rect 50300 68518 50346 68570
rect 50346 68518 50356 68570
rect 50380 68518 50410 68570
rect 50410 68518 50422 68570
rect 50422 68518 50436 68570
rect 50460 68518 50474 68570
rect 50474 68518 50486 68570
rect 50486 68518 50516 68570
rect 50540 68518 50550 68570
rect 50550 68518 50596 68570
rect 50300 68516 50356 68518
rect 50380 68516 50436 68518
rect 50460 68516 50516 68518
rect 50540 68516 50596 68518
rect 50300 67482 50356 67484
rect 50380 67482 50436 67484
rect 50460 67482 50516 67484
rect 50540 67482 50596 67484
rect 50300 67430 50346 67482
rect 50346 67430 50356 67482
rect 50380 67430 50410 67482
rect 50410 67430 50422 67482
rect 50422 67430 50436 67482
rect 50460 67430 50474 67482
rect 50474 67430 50486 67482
rect 50486 67430 50516 67482
rect 50540 67430 50550 67482
rect 50550 67430 50596 67482
rect 50300 67428 50356 67430
rect 50380 67428 50436 67430
rect 50460 67428 50516 67430
rect 50540 67428 50596 67430
rect 50300 66394 50356 66396
rect 50380 66394 50436 66396
rect 50460 66394 50516 66396
rect 50540 66394 50596 66396
rect 50300 66342 50346 66394
rect 50346 66342 50356 66394
rect 50380 66342 50410 66394
rect 50410 66342 50422 66394
rect 50422 66342 50436 66394
rect 50460 66342 50474 66394
rect 50474 66342 50486 66394
rect 50486 66342 50516 66394
rect 50540 66342 50550 66394
rect 50550 66342 50596 66394
rect 50300 66340 50356 66342
rect 50380 66340 50436 66342
rect 50460 66340 50516 66342
rect 50540 66340 50596 66342
rect 50300 65306 50356 65308
rect 50380 65306 50436 65308
rect 50460 65306 50516 65308
rect 50540 65306 50596 65308
rect 50300 65254 50346 65306
rect 50346 65254 50356 65306
rect 50380 65254 50410 65306
rect 50410 65254 50422 65306
rect 50422 65254 50436 65306
rect 50460 65254 50474 65306
rect 50474 65254 50486 65306
rect 50486 65254 50516 65306
rect 50540 65254 50550 65306
rect 50550 65254 50596 65306
rect 50300 65252 50356 65254
rect 50380 65252 50436 65254
rect 50460 65252 50516 65254
rect 50540 65252 50596 65254
rect 50300 64218 50356 64220
rect 50380 64218 50436 64220
rect 50460 64218 50516 64220
rect 50540 64218 50596 64220
rect 50300 64166 50346 64218
rect 50346 64166 50356 64218
rect 50380 64166 50410 64218
rect 50410 64166 50422 64218
rect 50422 64166 50436 64218
rect 50460 64166 50474 64218
rect 50474 64166 50486 64218
rect 50486 64166 50516 64218
rect 50540 64166 50550 64218
rect 50550 64166 50596 64218
rect 50300 64164 50356 64166
rect 50380 64164 50436 64166
rect 50460 64164 50516 64166
rect 50540 64164 50596 64166
rect 50300 63130 50356 63132
rect 50380 63130 50436 63132
rect 50460 63130 50516 63132
rect 50540 63130 50596 63132
rect 50300 63078 50346 63130
rect 50346 63078 50356 63130
rect 50380 63078 50410 63130
rect 50410 63078 50422 63130
rect 50422 63078 50436 63130
rect 50460 63078 50474 63130
rect 50474 63078 50486 63130
rect 50486 63078 50516 63130
rect 50540 63078 50550 63130
rect 50550 63078 50596 63130
rect 50300 63076 50356 63078
rect 50380 63076 50436 63078
rect 50460 63076 50516 63078
rect 50540 63076 50596 63078
rect 50300 62042 50356 62044
rect 50380 62042 50436 62044
rect 50460 62042 50516 62044
rect 50540 62042 50596 62044
rect 50300 61990 50346 62042
rect 50346 61990 50356 62042
rect 50380 61990 50410 62042
rect 50410 61990 50422 62042
rect 50422 61990 50436 62042
rect 50460 61990 50474 62042
rect 50474 61990 50486 62042
rect 50486 61990 50516 62042
rect 50540 61990 50550 62042
rect 50550 61990 50596 62042
rect 50300 61988 50356 61990
rect 50380 61988 50436 61990
rect 50460 61988 50516 61990
rect 50540 61988 50596 61990
rect 50300 60954 50356 60956
rect 50380 60954 50436 60956
rect 50460 60954 50516 60956
rect 50540 60954 50596 60956
rect 50300 60902 50346 60954
rect 50346 60902 50356 60954
rect 50380 60902 50410 60954
rect 50410 60902 50422 60954
rect 50422 60902 50436 60954
rect 50460 60902 50474 60954
rect 50474 60902 50486 60954
rect 50486 60902 50516 60954
rect 50540 60902 50550 60954
rect 50550 60902 50596 60954
rect 50300 60900 50356 60902
rect 50380 60900 50436 60902
rect 50460 60900 50516 60902
rect 50540 60900 50596 60902
rect 50300 59866 50356 59868
rect 50380 59866 50436 59868
rect 50460 59866 50516 59868
rect 50540 59866 50596 59868
rect 50300 59814 50346 59866
rect 50346 59814 50356 59866
rect 50380 59814 50410 59866
rect 50410 59814 50422 59866
rect 50422 59814 50436 59866
rect 50460 59814 50474 59866
rect 50474 59814 50486 59866
rect 50486 59814 50516 59866
rect 50540 59814 50550 59866
rect 50550 59814 50596 59866
rect 50300 59812 50356 59814
rect 50380 59812 50436 59814
rect 50460 59812 50516 59814
rect 50540 59812 50596 59814
rect 50300 58778 50356 58780
rect 50380 58778 50436 58780
rect 50460 58778 50516 58780
rect 50540 58778 50596 58780
rect 50300 58726 50346 58778
rect 50346 58726 50356 58778
rect 50380 58726 50410 58778
rect 50410 58726 50422 58778
rect 50422 58726 50436 58778
rect 50460 58726 50474 58778
rect 50474 58726 50486 58778
rect 50486 58726 50516 58778
rect 50540 58726 50550 58778
rect 50550 58726 50596 58778
rect 50300 58724 50356 58726
rect 50380 58724 50436 58726
rect 50460 58724 50516 58726
rect 50540 58724 50596 58726
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 2870 720 2926 776
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 65660 69114 65716 69116
rect 65740 69114 65796 69116
rect 65820 69114 65876 69116
rect 65900 69114 65956 69116
rect 65660 69062 65706 69114
rect 65706 69062 65716 69114
rect 65740 69062 65770 69114
rect 65770 69062 65782 69114
rect 65782 69062 65796 69114
rect 65820 69062 65834 69114
rect 65834 69062 65846 69114
rect 65846 69062 65876 69114
rect 65900 69062 65910 69114
rect 65910 69062 65956 69114
rect 65660 69060 65716 69062
rect 65740 69060 65796 69062
rect 65820 69060 65876 69062
rect 65900 69060 65956 69062
rect 65660 68026 65716 68028
rect 65740 68026 65796 68028
rect 65820 68026 65876 68028
rect 65900 68026 65956 68028
rect 65660 67974 65706 68026
rect 65706 67974 65716 68026
rect 65740 67974 65770 68026
rect 65770 67974 65782 68026
rect 65782 67974 65796 68026
rect 65820 67974 65834 68026
rect 65834 67974 65846 68026
rect 65846 67974 65876 68026
rect 65900 67974 65910 68026
rect 65910 67974 65956 68026
rect 65660 67972 65716 67974
rect 65740 67972 65796 67974
rect 65820 67972 65876 67974
rect 65900 67972 65956 67974
rect 67730 70080 67786 70136
rect 65660 66938 65716 66940
rect 65740 66938 65796 66940
rect 65820 66938 65876 66940
rect 65900 66938 65956 66940
rect 65660 66886 65706 66938
rect 65706 66886 65716 66938
rect 65740 66886 65770 66938
rect 65770 66886 65782 66938
rect 65782 66886 65796 66938
rect 65820 66886 65834 66938
rect 65834 66886 65846 66938
rect 65846 66886 65876 66938
rect 65900 66886 65910 66938
rect 65910 66886 65956 66938
rect 65660 66884 65716 66886
rect 65740 66884 65796 66886
rect 65820 66884 65876 66886
rect 65900 66884 65956 66886
rect 65660 65850 65716 65852
rect 65740 65850 65796 65852
rect 65820 65850 65876 65852
rect 65900 65850 65956 65852
rect 65660 65798 65706 65850
rect 65706 65798 65716 65850
rect 65740 65798 65770 65850
rect 65770 65798 65782 65850
rect 65782 65798 65796 65850
rect 65820 65798 65834 65850
rect 65834 65798 65846 65850
rect 65846 65798 65876 65850
rect 65900 65798 65910 65850
rect 65910 65798 65956 65850
rect 65660 65796 65716 65798
rect 65740 65796 65796 65798
rect 65820 65796 65876 65798
rect 65900 65796 65956 65798
rect 65660 64762 65716 64764
rect 65740 64762 65796 64764
rect 65820 64762 65876 64764
rect 65900 64762 65956 64764
rect 65660 64710 65706 64762
rect 65706 64710 65716 64762
rect 65740 64710 65770 64762
rect 65770 64710 65782 64762
rect 65782 64710 65796 64762
rect 65820 64710 65834 64762
rect 65834 64710 65846 64762
rect 65846 64710 65876 64762
rect 65900 64710 65910 64762
rect 65910 64710 65956 64762
rect 65660 64708 65716 64710
rect 65740 64708 65796 64710
rect 65820 64708 65876 64710
rect 65900 64708 65956 64710
rect 65660 63674 65716 63676
rect 65740 63674 65796 63676
rect 65820 63674 65876 63676
rect 65900 63674 65956 63676
rect 65660 63622 65706 63674
rect 65706 63622 65716 63674
rect 65740 63622 65770 63674
rect 65770 63622 65782 63674
rect 65782 63622 65796 63674
rect 65820 63622 65834 63674
rect 65834 63622 65846 63674
rect 65846 63622 65876 63674
rect 65900 63622 65910 63674
rect 65910 63622 65956 63674
rect 65660 63620 65716 63622
rect 65740 63620 65796 63622
rect 65820 63620 65876 63622
rect 65900 63620 65956 63622
rect 65660 62586 65716 62588
rect 65740 62586 65796 62588
rect 65820 62586 65876 62588
rect 65900 62586 65956 62588
rect 65660 62534 65706 62586
rect 65706 62534 65716 62586
rect 65740 62534 65770 62586
rect 65770 62534 65782 62586
rect 65782 62534 65796 62586
rect 65820 62534 65834 62586
rect 65834 62534 65846 62586
rect 65846 62534 65876 62586
rect 65900 62534 65910 62586
rect 65910 62534 65956 62586
rect 65660 62532 65716 62534
rect 65740 62532 65796 62534
rect 65820 62532 65876 62534
rect 65900 62532 65956 62534
rect 65660 61498 65716 61500
rect 65740 61498 65796 61500
rect 65820 61498 65876 61500
rect 65900 61498 65956 61500
rect 65660 61446 65706 61498
rect 65706 61446 65716 61498
rect 65740 61446 65770 61498
rect 65770 61446 65782 61498
rect 65782 61446 65796 61498
rect 65820 61446 65834 61498
rect 65834 61446 65846 61498
rect 65846 61446 65876 61498
rect 65900 61446 65910 61498
rect 65910 61446 65956 61498
rect 65660 61444 65716 61446
rect 65740 61444 65796 61446
rect 65820 61444 65876 61446
rect 65900 61444 65956 61446
rect 65660 60410 65716 60412
rect 65740 60410 65796 60412
rect 65820 60410 65876 60412
rect 65900 60410 65956 60412
rect 65660 60358 65706 60410
rect 65706 60358 65716 60410
rect 65740 60358 65770 60410
rect 65770 60358 65782 60410
rect 65782 60358 65796 60410
rect 65820 60358 65834 60410
rect 65834 60358 65846 60410
rect 65846 60358 65876 60410
rect 65900 60358 65910 60410
rect 65910 60358 65956 60410
rect 65660 60356 65716 60358
rect 65740 60356 65796 60358
rect 65820 60356 65876 60358
rect 65900 60356 65956 60358
rect 65660 59322 65716 59324
rect 65740 59322 65796 59324
rect 65820 59322 65876 59324
rect 65900 59322 65956 59324
rect 65660 59270 65706 59322
rect 65706 59270 65716 59322
rect 65740 59270 65770 59322
rect 65770 59270 65782 59322
rect 65782 59270 65796 59322
rect 65820 59270 65834 59322
rect 65834 59270 65846 59322
rect 65846 59270 65876 59322
rect 65900 59270 65910 59322
rect 65910 59270 65956 59322
rect 65660 59268 65716 59270
rect 65740 59268 65796 59270
rect 65820 59268 65876 59270
rect 65900 59268 65956 59270
rect 65660 58234 65716 58236
rect 65740 58234 65796 58236
rect 65820 58234 65876 58236
rect 65900 58234 65956 58236
rect 65660 58182 65706 58234
rect 65706 58182 65716 58234
rect 65740 58182 65770 58234
rect 65770 58182 65782 58234
rect 65782 58182 65796 58234
rect 65820 58182 65834 58234
rect 65834 58182 65846 58234
rect 65846 58182 65876 58234
rect 65900 58182 65910 58234
rect 65910 58182 65956 58234
rect 65660 58180 65716 58182
rect 65740 58180 65796 58182
rect 65820 58180 65876 58182
rect 65900 58180 65956 58182
rect 65660 57146 65716 57148
rect 65740 57146 65796 57148
rect 65820 57146 65876 57148
rect 65900 57146 65956 57148
rect 65660 57094 65706 57146
rect 65706 57094 65716 57146
rect 65740 57094 65770 57146
rect 65770 57094 65782 57146
rect 65782 57094 65796 57146
rect 65820 57094 65834 57146
rect 65834 57094 65846 57146
rect 65846 57094 65876 57146
rect 65900 57094 65910 57146
rect 65910 57094 65956 57146
rect 65660 57092 65716 57094
rect 65740 57092 65796 57094
rect 65820 57092 65876 57094
rect 65900 57092 65956 57094
rect 65660 56058 65716 56060
rect 65740 56058 65796 56060
rect 65820 56058 65876 56060
rect 65900 56058 65956 56060
rect 65660 56006 65706 56058
rect 65706 56006 65716 56058
rect 65740 56006 65770 56058
rect 65770 56006 65782 56058
rect 65782 56006 65796 56058
rect 65820 56006 65834 56058
rect 65834 56006 65846 56058
rect 65846 56006 65876 56058
rect 65900 56006 65910 56058
rect 65910 56006 65956 56058
rect 65660 56004 65716 56006
rect 65740 56004 65796 56006
rect 65820 56004 65876 56006
rect 65900 56004 65956 56006
rect 66166 55120 66222 55176
rect 65660 54970 65716 54972
rect 65740 54970 65796 54972
rect 65820 54970 65876 54972
rect 65900 54970 65956 54972
rect 65660 54918 65706 54970
rect 65706 54918 65716 54970
rect 65740 54918 65770 54970
rect 65770 54918 65782 54970
rect 65782 54918 65796 54970
rect 65820 54918 65834 54970
rect 65834 54918 65846 54970
rect 65846 54918 65876 54970
rect 65900 54918 65910 54970
rect 65910 54918 65956 54970
rect 65660 54916 65716 54918
rect 65740 54916 65796 54918
rect 65820 54916 65876 54918
rect 65900 54916 65956 54918
rect 65660 53882 65716 53884
rect 65740 53882 65796 53884
rect 65820 53882 65876 53884
rect 65900 53882 65956 53884
rect 65660 53830 65706 53882
rect 65706 53830 65716 53882
rect 65740 53830 65770 53882
rect 65770 53830 65782 53882
rect 65782 53830 65796 53882
rect 65820 53830 65834 53882
rect 65834 53830 65846 53882
rect 65846 53830 65876 53882
rect 65900 53830 65910 53882
rect 65910 53830 65956 53882
rect 65660 53828 65716 53830
rect 65740 53828 65796 53830
rect 65820 53828 65876 53830
rect 65900 53828 65956 53830
rect 65660 52794 65716 52796
rect 65740 52794 65796 52796
rect 65820 52794 65876 52796
rect 65900 52794 65956 52796
rect 65660 52742 65706 52794
rect 65706 52742 65716 52794
rect 65740 52742 65770 52794
rect 65770 52742 65782 52794
rect 65782 52742 65796 52794
rect 65820 52742 65834 52794
rect 65834 52742 65846 52794
rect 65846 52742 65876 52794
rect 65900 52742 65910 52794
rect 65910 52742 65956 52794
rect 65660 52740 65716 52742
rect 65740 52740 65796 52742
rect 65820 52740 65876 52742
rect 65900 52740 65956 52742
rect 65660 51706 65716 51708
rect 65740 51706 65796 51708
rect 65820 51706 65876 51708
rect 65900 51706 65956 51708
rect 65660 51654 65706 51706
rect 65706 51654 65716 51706
rect 65740 51654 65770 51706
rect 65770 51654 65782 51706
rect 65782 51654 65796 51706
rect 65820 51654 65834 51706
rect 65834 51654 65846 51706
rect 65846 51654 65876 51706
rect 65900 51654 65910 51706
rect 65910 51654 65956 51706
rect 65660 51652 65716 51654
rect 65740 51652 65796 51654
rect 65820 51652 65876 51654
rect 65900 51652 65956 51654
rect 65660 50618 65716 50620
rect 65740 50618 65796 50620
rect 65820 50618 65876 50620
rect 65900 50618 65956 50620
rect 65660 50566 65706 50618
rect 65706 50566 65716 50618
rect 65740 50566 65770 50618
rect 65770 50566 65782 50618
rect 65782 50566 65796 50618
rect 65820 50566 65834 50618
rect 65834 50566 65846 50618
rect 65846 50566 65876 50618
rect 65900 50566 65910 50618
rect 65910 50566 65956 50618
rect 65660 50564 65716 50566
rect 65740 50564 65796 50566
rect 65820 50564 65876 50566
rect 65900 50564 65956 50566
rect 65522 49680 65578 49736
rect 65660 49530 65716 49532
rect 65740 49530 65796 49532
rect 65820 49530 65876 49532
rect 65900 49530 65956 49532
rect 65660 49478 65706 49530
rect 65706 49478 65716 49530
rect 65740 49478 65770 49530
rect 65770 49478 65782 49530
rect 65782 49478 65796 49530
rect 65820 49478 65834 49530
rect 65834 49478 65846 49530
rect 65846 49478 65876 49530
rect 65900 49478 65910 49530
rect 65910 49478 65956 49530
rect 65660 49476 65716 49478
rect 65740 49476 65796 49478
rect 65820 49476 65876 49478
rect 65900 49476 65956 49478
rect 65660 48442 65716 48444
rect 65740 48442 65796 48444
rect 65820 48442 65876 48444
rect 65900 48442 65956 48444
rect 65660 48390 65706 48442
rect 65706 48390 65716 48442
rect 65740 48390 65770 48442
rect 65770 48390 65782 48442
rect 65782 48390 65796 48442
rect 65820 48390 65834 48442
rect 65834 48390 65846 48442
rect 65846 48390 65876 48442
rect 65900 48390 65910 48442
rect 65910 48390 65956 48442
rect 65660 48388 65716 48390
rect 65740 48388 65796 48390
rect 65820 48388 65876 48390
rect 65900 48388 65956 48390
rect 65660 47354 65716 47356
rect 65740 47354 65796 47356
rect 65820 47354 65876 47356
rect 65900 47354 65956 47356
rect 65660 47302 65706 47354
rect 65706 47302 65716 47354
rect 65740 47302 65770 47354
rect 65770 47302 65782 47354
rect 65782 47302 65796 47354
rect 65820 47302 65834 47354
rect 65834 47302 65846 47354
rect 65846 47302 65876 47354
rect 65900 47302 65910 47354
rect 65910 47302 65956 47354
rect 65660 47300 65716 47302
rect 65740 47300 65796 47302
rect 65820 47300 65876 47302
rect 65900 47300 65956 47302
rect 65660 46266 65716 46268
rect 65740 46266 65796 46268
rect 65820 46266 65876 46268
rect 65900 46266 65956 46268
rect 65660 46214 65706 46266
rect 65706 46214 65716 46266
rect 65740 46214 65770 46266
rect 65770 46214 65782 46266
rect 65782 46214 65796 46266
rect 65820 46214 65834 46266
rect 65834 46214 65846 46266
rect 65846 46214 65876 46266
rect 65900 46214 65910 46266
rect 65910 46214 65956 46266
rect 65660 46212 65716 46214
rect 65740 46212 65796 46214
rect 65820 46212 65876 46214
rect 65900 46212 65956 46214
rect 65660 45178 65716 45180
rect 65740 45178 65796 45180
rect 65820 45178 65876 45180
rect 65900 45178 65956 45180
rect 65660 45126 65706 45178
rect 65706 45126 65716 45178
rect 65740 45126 65770 45178
rect 65770 45126 65782 45178
rect 65782 45126 65796 45178
rect 65820 45126 65834 45178
rect 65834 45126 65846 45178
rect 65846 45126 65876 45178
rect 65900 45126 65910 45178
rect 65910 45126 65956 45178
rect 65660 45124 65716 45126
rect 65740 45124 65796 45126
rect 65820 45124 65876 45126
rect 65900 45124 65956 45126
rect 65660 44090 65716 44092
rect 65740 44090 65796 44092
rect 65820 44090 65876 44092
rect 65900 44090 65956 44092
rect 65660 44038 65706 44090
rect 65706 44038 65716 44090
rect 65740 44038 65770 44090
rect 65770 44038 65782 44090
rect 65782 44038 65796 44090
rect 65820 44038 65834 44090
rect 65834 44038 65846 44090
rect 65846 44038 65876 44090
rect 65900 44038 65910 44090
rect 65910 44038 65956 44090
rect 65660 44036 65716 44038
rect 65740 44036 65796 44038
rect 65820 44036 65876 44038
rect 65900 44036 65956 44038
rect 65660 43002 65716 43004
rect 65740 43002 65796 43004
rect 65820 43002 65876 43004
rect 65900 43002 65956 43004
rect 65660 42950 65706 43002
rect 65706 42950 65716 43002
rect 65740 42950 65770 43002
rect 65770 42950 65782 43002
rect 65782 42950 65796 43002
rect 65820 42950 65834 43002
rect 65834 42950 65846 43002
rect 65846 42950 65876 43002
rect 65900 42950 65910 43002
rect 65910 42950 65956 43002
rect 65660 42948 65716 42950
rect 65740 42948 65796 42950
rect 65820 42948 65876 42950
rect 65900 42948 65956 42950
rect 65660 41914 65716 41916
rect 65740 41914 65796 41916
rect 65820 41914 65876 41916
rect 65900 41914 65956 41916
rect 65660 41862 65706 41914
rect 65706 41862 65716 41914
rect 65740 41862 65770 41914
rect 65770 41862 65782 41914
rect 65782 41862 65796 41914
rect 65820 41862 65834 41914
rect 65834 41862 65846 41914
rect 65846 41862 65876 41914
rect 65900 41862 65910 41914
rect 65910 41862 65956 41914
rect 65660 41860 65716 41862
rect 65740 41860 65796 41862
rect 65820 41860 65876 41862
rect 65900 41860 65956 41862
rect 65660 40826 65716 40828
rect 65740 40826 65796 40828
rect 65820 40826 65876 40828
rect 65900 40826 65956 40828
rect 65660 40774 65706 40826
rect 65706 40774 65716 40826
rect 65740 40774 65770 40826
rect 65770 40774 65782 40826
rect 65782 40774 65796 40826
rect 65820 40774 65834 40826
rect 65834 40774 65846 40826
rect 65846 40774 65876 40826
rect 65900 40774 65910 40826
rect 65910 40774 65956 40826
rect 65660 40772 65716 40774
rect 65740 40772 65796 40774
rect 65820 40772 65876 40774
rect 65900 40772 65956 40774
rect 65660 39738 65716 39740
rect 65740 39738 65796 39740
rect 65820 39738 65876 39740
rect 65900 39738 65956 39740
rect 65660 39686 65706 39738
rect 65706 39686 65716 39738
rect 65740 39686 65770 39738
rect 65770 39686 65782 39738
rect 65782 39686 65796 39738
rect 65820 39686 65834 39738
rect 65834 39686 65846 39738
rect 65846 39686 65876 39738
rect 65900 39686 65910 39738
rect 65910 39686 65956 39738
rect 65660 39684 65716 39686
rect 65740 39684 65796 39686
rect 65820 39684 65876 39686
rect 65900 39684 65956 39686
rect 65660 38650 65716 38652
rect 65740 38650 65796 38652
rect 65820 38650 65876 38652
rect 65900 38650 65956 38652
rect 65660 38598 65706 38650
rect 65706 38598 65716 38650
rect 65740 38598 65770 38650
rect 65770 38598 65782 38650
rect 65782 38598 65796 38650
rect 65820 38598 65834 38650
rect 65834 38598 65846 38650
rect 65846 38598 65876 38650
rect 65900 38598 65910 38650
rect 65910 38598 65956 38650
rect 65660 38596 65716 38598
rect 65740 38596 65796 38598
rect 65820 38596 65876 38598
rect 65900 38596 65956 38598
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 66166 29960 66222 30016
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 67638 67360 67694 67416
rect 67270 59200 67326 59256
rect 67270 39480 67326 39536
rect 67546 66036 67548 66056
rect 67548 66036 67600 66056
rect 67600 66036 67602 66056
rect 67546 66000 67602 66036
rect 68098 63316 68100 63336
rect 68100 63316 68152 63336
rect 68152 63316 68154 63336
rect 68098 63280 68154 63316
rect 67638 61920 67694 61976
rect 67546 60596 67548 60616
rect 67548 60596 67600 60616
rect 67600 60596 67602 60616
rect 67546 60560 67602 60596
rect 68098 57876 68100 57896
rect 68100 57876 68152 57896
rect 68152 57876 68154 57896
rect 68098 57840 68154 57876
rect 67546 56480 67602 56536
rect 68098 51040 68154 51096
rect 67730 47640 67786 47696
rect 67546 46280 67602 46336
rect 68098 44940 68154 44976
rect 68098 44920 68100 44940
rect 68100 44920 68152 44940
rect 68152 44920 68154 44940
rect 68098 43560 68154 43616
rect 67546 42200 67602 42256
rect 68098 40840 68154 40896
rect 67546 35400 67602 35456
rect 67270 34040 67326 34096
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 66166 15680 66222 15736
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 68098 32680 68154 32736
rect 67546 31320 67602 31376
rect 68098 23180 68154 23216
rect 68098 23160 68100 23180
rect 68100 23160 68152 23180
rect 68152 23160 68154 23180
rect 67546 21120 67602 21176
rect 67822 18400 67878 18456
rect 67546 17076 67548 17096
rect 67548 17076 67600 17096
rect 67600 17076 67602 17096
rect 67546 17040 67602 17076
rect 67546 14320 67602 14376
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 67822 12960 67878 13016
rect 67638 7520 67694 7576
rect 67546 6196 67548 6216
rect 67548 6196 67600 6216
rect 67600 6196 67602 6216
rect 67546 6160 67602 6196
rect 67546 4800 67602 4856
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 66166 720 66222 776
<< metal3 >>
rect 0 71498 800 71588
rect 0 71348 858 71498
rect 69200 71348 70000 71588
rect 614 71302 858 71348
rect 614 70954 674 71302
rect 1393 70954 1459 70957
rect 614 70952 1459 70954
rect 614 70896 1398 70952
rect 1454 70896 1459 70952
rect 614 70894 1459 70896
rect 1393 70891 1459 70894
rect 0 69988 800 70228
rect 67725 70138 67791 70141
rect 69200 70138 70000 70228
rect 67725 70136 70000 70138
rect 67725 70080 67730 70136
rect 67786 70080 70000 70136
rect 67725 70078 70000 70080
rect 67725 70075 67791 70078
rect 69200 69988 70000 70078
rect 19568 69664 19888 69665
rect 19568 69600 19576 69664
rect 19640 69600 19656 69664
rect 19720 69600 19736 69664
rect 19800 69600 19816 69664
rect 19880 69600 19888 69664
rect 19568 69599 19888 69600
rect 50288 69664 50608 69665
rect 50288 69600 50296 69664
rect 50360 69600 50376 69664
rect 50440 69600 50456 69664
rect 50520 69600 50536 69664
rect 50600 69600 50608 69664
rect 50288 69599 50608 69600
rect 4208 69120 4528 69121
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 69055 4528 69056
rect 34928 69120 35248 69121
rect 34928 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35248 69120
rect 34928 69055 35248 69056
rect 65648 69120 65968 69121
rect 65648 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65968 69120
rect 65648 69055 65968 69056
rect 0 68778 800 68868
rect 2773 68778 2839 68781
rect 0 68776 2839 68778
rect 0 68720 2778 68776
rect 2834 68720 2839 68776
rect 0 68718 2839 68720
rect 0 68628 800 68718
rect 2773 68715 2839 68718
rect 69200 68628 70000 68868
rect 19568 68576 19888 68577
rect 19568 68512 19576 68576
rect 19640 68512 19656 68576
rect 19720 68512 19736 68576
rect 19800 68512 19816 68576
rect 19880 68512 19888 68576
rect 19568 68511 19888 68512
rect 50288 68576 50608 68577
rect 50288 68512 50296 68576
rect 50360 68512 50376 68576
rect 50440 68512 50456 68576
rect 50520 68512 50536 68576
rect 50600 68512 50608 68576
rect 50288 68511 50608 68512
rect 4208 68032 4528 68033
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 67967 4528 67968
rect 34928 68032 35248 68033
rect 34928 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35248 68032
rect 34928 67967 35248 67968
rect 65648 68032 65968 68033
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 67967 65968 67968
rect 0 67418 800 67508
rect 19568 67488 19888 67489
rect 19568 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19888 67488
rect 19568 67423 19888 67424
rect 50288 67488 50608 67489
rect 50288 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50608 67488
rect 50288 67423 50608 67424
rect 2773 67418 2839 67421
rect 0 67416 2839 67418
rect 0 67360 2778 67416
rect 2834 67360 2839 67416
rect 0 67358 2839 67360
rect 0 67268 800 67358
rect 2773 67355 2839 67358
rect 67633 67418 67699 67421
rect 69200 67418 70000 67508
rect 67633 67416 70000 67418
rect 67633 67360 67638 67416
rect 67694 67360 70000 67416
rect 67633 67358 70000 67360
rect 67633 67355 67699 67358
rect 69200 67268 70000 67358
rect 4208 66944 4528 66945
rect 4208 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4528 66944
rect 4208 66879 4528 66880
rect 34928 66944 35248 66945
rect 34928 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35248 66944
rect 34928 66879 35248 66880
rect 65648 66944 65968 66945
rect 65648 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65968 66944
rect 65648 66879 65968 66880
rect 19568 66400 19888 66401
rect 19568 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19888 66400
rect 19568 66335 19888 66336
rect 50288 66400 50608 66401
rect 50288 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50608 66400
rect 50288 66335 50608 66336
rect 0 65908 800 66148
rect 67541 66058 67607 66061
rect 69200 66058 70000 66148
rect 67541 66056 70000 66058
rect 67541 66000 67546 66056
rect 67602 66000 70000 66056
rect 67541 65998 70000 66000
rect 67541 65995 67607 65998
rect 69200 65908 70000 65998
rect 4208 65856 4528 65857
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 65791 4528 65792
rect 34928 65856 35248 65857
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 65791 35248 65792
rect 65648 65856 65968 65857
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 65791 65968 65792
rect 19568 65312 19888 65313
rect 19568 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19888 65312
rect 19568 65247 19888 65248
rect 50288 65312 50608 65313
rect 50288 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50608 65312
rect 50288 65247 50608 65248
rect 0 64548 800 64788
rect 4208 64768 4528 64769
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 64703 4528 64704
rect 34928 64768 35248 64769
rect 34928 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35248 64768
rect 34928 64703 35248 64704
rect 65648 64768 65968 64769
rect 65648 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65968 64768
rect 65648 64703 65968 64704
rect 69200 64548 70000 64788
rect 19568 64224 19888 64225
rect 19568 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19888 64224
rect 19568 64159 19888 64160
rect 50288 64224 50608 64225
rect 50288 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50608 64224
rect 50288 64159 50608 64160
rect 4208 63680 4528 63681
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 63615 4528 63616
rect 34928 63680 35248 63681
rect 34928 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35248 63680
rect 34928 63615 35248 63616
rect 65648 63680 65968 63681
rect 65648 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65968 63680
rect 65648 63615 65968 63616
rect 0 63338 800 63428
rect 1393 63338 1459 63341
rect 0 63336 1459 63338
rect 0 63280 1398 63336
rect 1454 63280 1459 63336
rect 0 63278 1459 63280
rect 0 63188 800 63278
rect 1393 63275 1459 63278
rect 68093 63338 68159 63341
rect 69200 63338 70000 63428
rect 68093 63336 70000 63338
rect 68093 63280 68098 63336
rect 68154 63280 70000 63336
rect 68093 63278 70000 63280
rect 68093 63275 68159 63278
rect 69200 63188 70000 63278
rect 19568 63136 19888 63137
rect 19568 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19888 63136
rect 19568 63071 19888 63072
rect 50288 63136 50608 63137
rect 50288 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50608 63136
rect 50288 63071 50608 63072
rect 4208 62592 4528 62593
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 62527 4528 62528
rect 34928 62592 35248 62593
rect 34928 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35248 62592
rect 34928 62527 35248 62528
rect 65648 62592 65968 62593
rect 65648 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65968 62592
rect 65648 62527 65968 62528
rect 0 61828 800 62068
rect 19568 62048 19888 62049
rect 19568 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19888 62048
rect 19568 61983 19888 61984
rect 50288 62048 50608 62049
rect 50288 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50608 62048
rect 50288 61983 50608 61984
rect 67633 61978 67699 61981
rect 69200 61978 70000 62068
rect 67633 61976 70000 61978
rect 67633 61920 67638 61976
rect 67694 61920 70000 61976
rect 67633 61918 70000 61920
rect 67633 61915 67699 61918
rect 69200 61828 70000 61918
rect 4208 61504 4528 61505
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 61439 4528 61440
rect 34928 61504 35248 61505
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 34928 61439 35248 61440
rect 65648 61504 65968 61505
rect 65648 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65968 61504
rect 65648 61439 65968 61440
rect 19568 60960 19888 60961
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 60895 19888 60896
rect 50288 60960 50608 60961
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 60895 50608 60896
rect 0 60618 800 60708
rect 1853 60618 1919 60621
rect 0 60616 1919 60618
rect 0 60560 1858 60616
rect 1914 60560 1919 60616
rect 0 60558 1919 60560
rect 0 60468 800 60558
rect 1853 60555 1919 60558
rect 67541 60618 67607 60621
rect 69200 60618 70000 60708
rect 67541 60616 70000 60618
rect 67541 60560 67546 60616
rect 67602 60560 70000 60616
rect 67541 60558 70000 60560
rect 67541 60555 67607 60558
rect 69200 60468 70000 60558
rect 4208 60416 4528 60417
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 60351 4528 60352
rect 34928 60416 35248 60417
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 60351 35248 60352
rect 65648 60416 65968 60417
rect 65648 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65968 60416
rect 65648 60351 65968 60352
rect 19568 59872 19888 59873
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 59807 19888 59808
rect 50288 59872 50608 59873
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 59807 50608 59808
rect 0 59258 800 59348
rect 4208 59328 4528 59329
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 59263 4528 59264
rect 34928 59328 35248 59329
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 59263 35248 59264
rect 65648 59328 65968 59329
rect 65648 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65968 59328
rect 65648 59263 65968 59264
rect 2773 59258 2839 59261
rect 0 59256 2839 59258
rect 0 59200 2778 59256
rect 2834 59200 2839 59256
rect 0 59198 2839 59200
rect 0 59108 800 59198
rect 2773 59195 2839 59198
rect 67265 59258 67331 59261
rect 69200 59258 70000 59348
rect 67265 59256 70000 59258
rect 67265 59200 67270 59256
rect 67326 59200 70000 59256
rect 67265 59198 70000 59200
rect 67265 59195 67331 59198
rect 69200 59108 70000 59198
rect 19568 58784 19888 58785
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 58719 19888 58720
rect 50288 58784 50608 58785
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 58719 50608 58720
rect 4208 58240 4528 58241
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 58175 4528 58176
rect 34928 58240 35248 58241
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 58175 35248 58176
rect 65648 58240 65968 58241
rect 65648 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65968 58240
rect 65648 58175 65968 58176
rect 0 57748 800 57988
rect 25998 57972 26004 58036
rect 26068 58034 26074 58036
rect 26141 58034 26207 58037
rect 26068 58032 26207 58034
rect 26068 57976 26146 58032
rect 26202 57976 26207 58032
rect 26068 57974 26207 57976
rect 26068 57972 26074 57974
rect 26141 57971 26207 57974
rect 68093 57898 68159 57901
rect 69200 57898 70000 57988
rect 68093 57896 70000 57898
rect 68093 57840 68098 57896
rect 68154 57840 70000 57896
rect 68093 57838 70000 57840
rect 68093 57835 68159 57838
rect 69200 57748 70000 57838
rect 19568 57696 19888 57697
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 57631 19888 57632
rect 50288 57696 50608 57697
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 57631 50608 57632
rect 4208 57152 4528 57153
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 57087 4528 57088
rect 34928 57152 35248 57153
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 57087 35248 57088
rect 65648 57152 65968 57153
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 57087 65968 57088
rect 0 56538 800 56628
rect 19568 56608 19888 56609
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 56543 19888 56544
rect 50288 56608 50608 56609
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 56543 50608 56544
rect 1393 56538 1459 56541
rect 0 56536 1459 56538
rect 0 56480 1398 56536
rect 1454 56480 1459 56536
rect 0 56478 1459 56480
rect 0 56388 800 56478
rect 1393 56475 1459 56478
rect 67541 56538 67607 56541
rect 69200 56538 70000 56628
rect 67541 56536 70000 56538
rect 67541 56480 67546 56536
rect 67602 56480 70000 56536
rect 67541 56478 70000 56480
rect 67541 56475 67607 56478
rect 69200 56388 70000 56478
rect 4208 56064 4528 56065
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 55999 4528 56000
rect 34928 56064 35248 56065
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 55999 35248 56000
rect 65648 56064 65968 56065
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 55999 65968 56000
rect 19568 55520 19888 55521
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 55455 19888 55456
rect 50288 55520 50608 55521
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 55455 50608 55456
rect 0 55178 800 55268
rect 3509 55178 3575 55181
rect 0 55176 3575 55178
rect 0 55120 3514 55176
rect 3570 55120 3575 55176
rect 0 55118 3575 55120
rect 0 55028 800 55118
rect 3509 55115 3575 55118
rect 66161 55178 66227 55181
rect 69200 55178 70000 55268
rect 66161 55176 70000 55178
rect 66161 55120 66166 55176
rect 66222 55120 70000 55176
rect 66161 55118 70000 55120
rect 66161 55115 66227 55118
rect 69200 55028 70000 55118
rect 4208 54976 4528 54977
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 54911 4528 54912
rect 34928 54976 35248 54977
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 54911 35248 54912
rect 65648 54976 65968 54977
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 54911 65968 54912
rect 19568 54432 19888 54433
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 54367 19888 54368
rect 50288 54432 50608 54433
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 54367 50608 54368
rect 0 53818 800 53908
rect 4208 53888 4528 53889
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 53823 4528 53824
rect 34928 53888 35248 53889
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 53823 35248 53824
rect 65648 53888 65968 53889
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 53823 65968 53824
rect 2773 53818 2839 53821
rect 0 53816 2839 53818
rect 0 53760 2778 53816
rect 2834 53760 2839 53816
rect 0 53758 2839 53760
rect 0 53668 800 53758
rect 2773 53755 2839 53758
rect 69200 53668 70000 53908
rect 19568 53344 19888 53345
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 53279 19888 53280
rect 50288 53344 50608 53345
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 53279 50608 53280
rect 41413 53002 41479 53005
rect 42701 53002 42767 53005
rect 41413 53000 42767 53002
rect 41413 52944 41418 53000
rect 41474 52944 42706 53000
rect 42762 52944 42767 53000
rect 41413 52942 42767 52944
rect 41413 52939 41479 52942
rect 42701 52939 42767 52942
rect 4208 52800 4528 52801
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 52735 4528 52736
rect 34928 52800 35248 52801
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 52735 35248 52736
rect 65648 52800 65968 52801
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 52735 65968 52736
rect 0 52458 800 52548
rect 1853 52458 1919 52461
rect 0 52456 1919 52458
rect 0 52400 1858 52456
rect 1914 52400 1919 52456
rect 0 52398 1919 52400
rect 0 52308 800 52398
rect 1853 52395 1919 52398
rect 69200 52308 70000 52548
rect 19568 52256 19888 52257
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 52191 19888 52192
rect 50288 52256 50608 52257
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 52191 50608 52192
rect 4208 51712 4528 51713
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 51647 4528 51648
rect 34928 51712 35248 51713
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 51647 35248 51648
rect 65648 51712 65968 51713
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 51647 65968 51648
rect 0 51098 800 51188
rect 19568 51168 19888 51169
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 51103 19888 51104
rect 50288 51168 50608 51169
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 51103 50608 51104
rect 3509 51098 3575 51101
rect 0 51096 3575 51098
rect 0 51040 3514 51096
rect 3570 51040 3575 51096
rect 0 51038 3575 51040
rect 0 50948 800 51038
rect 3509 51035 3575 51038
rect 68093 51098 68159 51101
rect 69200 51098 70000 51188
rect 68093 51096 70000 51098
rect 68093 51040 68098 51096
rect 68154 51040 70000 51096
rect 68093 51038 70000 51040
rect 68093 51035 68159 51038
rect 42609 50962 42675 50965
rect 43897 50962 43963 50965
rect 42609 50960 43963 50962
rect 42609 50904 42614 50960
rect 42670 50904 43902 50960
rect 43958 50904 43963 50960
rect 69200 50948 70000 51038
rect 42609 50902 43963 50904
rect 42609 50899 42675 50902
rect 43897 50899 43963 50902
rect 4208 50624 4528 50625
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 50559 4528 50560
rect 34928 50624 35248 50625
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 50559 35248 50560
rect 65648 50624 65968 50625
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 50559 65968 50560
rect 19568 50080 19888 50081
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 50015 19888 50016
rect 50288 50080 50608 50081
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 50015 50608 50016
rect 0 49738 800 49828
rect 3509 49738 3575 49741
rect 25865 49740 25931 49741
rect 25814 49738 25820 49740
rect 0 49736 3575 49738
rect 0 49680 3514 49736
rect 3570 49680 3575 49736
rect 0 49678 3575 49680
rect 25774 49678 25820 49738
rect 25884 49736 25931 49740
rect 25926 49680 25931 49736
rect 0 49588 800 49678
rect 3509 49675 3575 49678
rect 25814 49676 25820 49678
rect 25884 49676 25931 49680
rect 25865 49675 25931 49676
rect 65517 49738 65583 49741
rect 69200 49738 70000 49828
rect 65517 49736 70000 49738
rect 65517 49680 65522 49736
rect 65578 49680 70000 49736
rect 65517 49678 70000 49680
rect 65517 49675 65583 49678
rect 69200 49588 70000 49678
rect 4208 49536 4528 49537
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 49471 4528 49472
rect 34928 49536 35248 49537
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 49471 35248 49472
rect 65648 49536 65968 49537
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 49471 65968 49472
rect 34605 49330 34671 49333
rect 34881 49330 34947 49333
rect 34605 49328 34947 49330
rect 34605 49272 34610 49328
rect 34666 49272 34886 49328
rect 34942 49272 34947 49328
rect 34605 49270 34947 49272
rect 34605 49267 34671 49270
rect 34881 49267 34947 49270
rect 43713 49194 43779 49197
rect 45645 49194 45711 49197
rect 43713 49192 45711 49194
rect 43713 49136 43718 49192
rect 43774 49136 45650 49192
rect 45706 49136 45711 49192
rect 43713 49134 45711 49136
rect 43713 49131 43779 49134
rect 45645 49131 45711 49134
rect 19568 48992 19888 48993
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 48927 19888 48928
rect 50288 48992 50608 48993
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 48927 50608 48928
rect 0 48228 800 48468
rect 4208 48448 4528 48449
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 48383 4528 48384
rect 34928 48448 35248 48449
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 48383 35248 48384
rect 65648 48448 65968 48449
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 48383 65968 48384
rect 32949 48242 33015 48245
rect 33961 48242 34027 48245
rect 32949 48240 34027 48242
rect 32949 48184 32954 48240
rect 33010 48184 33966 48240
rect 34022 48184 34027 48240
rect 69200 48228 70000 48468
rect 32949 48182 34027 48184
rect 32949 48179 33015 48182
rect 33961 48179 34027 48182
rect 30281 48106 30347 48109
rect 36353 48106 36419 48109
rect 30281 48104 36419 48106
rect 30281 48048 30286 48104
rect 30342 48048 36358 48104
rect 36414 48048 36419 48104
rect 30281 48046 36419 48048
rect 30281 48043 30347 48046
rect 36353 48043 36419 48046
rect 33225 47970 33291 47973
rect 33869 47970 33935 47973
rect 33225 47968 33935 47970
rect 33225 47912 33230 47968
rect 33286 47912 33874 47968
rect 33930 47912 33935 47968
rect 33225 47910 33935 47912
rect 33225 47907 33291 47910
rect 33869 47907 33935 47910
rect 19568 47904 19888 47905
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 47839 19888 47840
rect 50288 47904 50608 47905
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 47839 50608 47840
rect 33777 47834 33843 47837
rect 35985 47834 36051 47837
rect 33777 47832 36051 47834
rect 0 47698 800 47788
rect 33777 47776 33782 47832
rect 33838 47776 35990 47832
rect 36046 47776 36051 47832
rect 33777 47774 36051 47776
rect 33777 47771 33843 47774
rect 35985 47771 36051 47774
rect 2773 47698 2839 47701
rect 0 47696 2839 47698
rect 0 47640 2778 47696
rect 2834 47640 2839 47696
rect 0 47638 2839 47640
rect 0 47548 800 47638
rect 2773 47635 2839 47638
rect 67725 47698 67791 47701
rect 69200 47698 70000 47788
rect 67725 47696 70000 47698
rect 67725 47640 67730 47696
rect 67786 47640 70000 47696
rect 67725 47638 70000 47640
rect 67725 47635 67791 47638
rect 69200 47548 70000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 65648 47360 65968 47361
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 47295 65968 47296
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 50288 46816 50608 46817
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 46751 50608 46752
rect 26049 46474 26115 46477
rect 26325 46474 26391 46477
rect 26049 46472 26391 46474
rect 0 46338 800 46428
rect 26049 46416 26054 46472
rect 26110 46416 26330 46472
rect 26386 46416 26391 46472
rect 26049 46414 26391 46416
rect 26049 46411 26115 46414
rect 26325 46411 26391 46414
rect 1853 46338 1919 46341
rect 0 46336 1919 46338
rect 0 46280 1858 46336
rect 1914 46280 1919 46336
rect 0 46278 1919 46280
rect 0 46188 800 46278
rect 1853 46275 1919 46278
rect 67541 46338 67607 46341
rect 69200 46338 70000 46428
rect 67541 46336 70000 46338
rect 67541 46280 67546 46336
rect 67602 46280 70000 46336
rect 67541 46278 70000 46280
rect 67541 46275 67607 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 65648 46272 65968 46273
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 46207 65968 46208
rect 69200 46188 70000 46278
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 50288 45728 50608 45729
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 45663 50608 45664
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 65648 45184 65968 45185
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 45119 65968 45120
rect 0 44978 800 45068
rect 1853 44978 1919 44981
rect 0 44976 1919 44978
rect 0 44920 1858 44976
rect 1914 44920 1919 44976
rect 0 44918 1919 44920
rect 0 44828 800 44918
rect 1853 44915 1919 44918
rect 68093 44978 68159 44981
rect 69200 44978 70000 45068
rect 68093 44976 70000 44978
rect 68093 44920 68098 44976
rect 68154 44920 70000 44976
rect 68093 44918 70000 44920
rect 68093 44915 68159 44918
rect 69200 44828 70000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 50288 44640 50608 44641
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 44575 50608 44576
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 65648 44096 65968 44097
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 44031 65968 44032
rect 0 43618 800 43708
rect 1853 43618 1919 43621
rect 0 43616 1919 43618
rect 0 43560 1858 43616
rect 1914 43560 1919 43616
rect 0 43558 1919 43560
rect 0 43468 800 43558
rect 1853 43555 1919 43558
rect 68093 43618 68159 43621
rect 69200 43618 70000 43708
rect 68093 43616 70000 43618
rect 68093 43560 68098 43616
rect 68154 43560 70000 43616
rect 68093 43558 70000 43560
rect 68093 43555 68159 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 50288 43552 50608 43553
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 43487 50608 43488
rect 69200 43468 70000 43558
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 65648 43008 65968 43009
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 42943 65968 42944
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 50288 42464 50608 42465
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 42399 50608 42400
rect 0 42258 800 42348
rect 1853 42258 1919 42261
rect 0 42256 1919 42258
rect 0 42200 1858 42256
rect 1914 42200 1919 42256
rect 0 42198 1919 42200
rect 0 42108 800 42198
rect 1853 42195 1919 42198
rect 2037 42258 2103 42261
rect 26141 42258 26207 42261
rect 2037 42256 26207 42258
rect 2037 42200 2042 42256
rect 2098 42200 26146 42256
rect 26202 42200 26207 42256
rect 2037 42198 26207 42200
rect 2037 42195 2103 42198
rect 26141 42195 26207 42198
rect 67541 42258 67607 42261
rect 69200 42258 70000 42348
rect 67541 42256 70000 42258
rect 67541 42200 67546 42256
rect 67602 42200 70000 42256
rect 67541 42198 70000 42200
rect 67541 42195 67607 42198
rect 69200 42108 70000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 65648 41920 65968 41921
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 41855 65968 41856
rect 37641 41850 37707 41853
rect 42241 41850 42307 41853
rect 37641 41848 42307 41850
rect 37641 41792 37646 41848
rect 37702 41792 42246 41848
rect 42302 41792 42307 41848
rect 37641 41790 42307 41792
rect 37641 41787 37707 41790
rect 42241 41787 42307 41790
rect 37273 41714 37339 41717
rect 39021 41714 39087 41717
rect 37273 41712 39087 41714
rect 37273 41656 37278 41712
rect 37334 41656 39026 41712
rect 39082 41656 39087 41712
rect 37273 41654 39087 41656
rect 37273 41651 37339 41654
rect 39021 41651 39087 41654
rect 21173 41578 21239 41581
rect 22461 41578 22527 41581
rect 28165 41578 28231 41581
rect 38101 41578 38167 41581
rect 21173 41576 28231 41578
rect 21173 41520 21178 41576
rect 21234 41520 22466 41576
rect 22522 41520 28170 41576
rect 28226 41520 28231 41576
rect 21173 41518 28231 41520
rect 21173 41515 21239 41518
rect 22461 41515 22527 41518
rect 28165 41515 28231 41518
rect 37782 41576 38167 41578
rect 37782 41520 38106 41576
rect 38162 41520 38167 41576
rect 37782 41518 38167 41520
rect 37641 41442 37707 41445
rect 37782 41442 37842 41518
rect 38101 41515 38167 41518
rect 37641 41440 37842 41442
rect 37641 41384 37646 41440
rect 37702 41384 37842 41440
rect 37641 41382 37842 41384
rect 37641 41379 37707 41382
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 50288 41376 50608 41377
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 41311 50608 41312
rect 38653 41170 38719 41173
rect 38653 41168 38762 41170
rect 38653 41112 38658 41168
rect 38714 41112 38762 41168
rect 38653 41107 38762 41112
rect 38702 41034 38762 41107
rect 40309 41034 40375 41037
rect 46381 41034 46447 41037
rect 38702 41032 46447 41034
rect 0 40898 800 40988
rect 38702 40976 40314 41032
rect 40370 40976 46386 41032
rect 46442 40976 46447 41032
rect 38702 40974 46447 40976
rect 40309 40971 40375 40974
rect 46381 40971 46447 40974
rect 3233 40898 3299 40901
rect 0 40896 3299 40898
rect 0 40840 3238 40896
rect 3294 40840 3299 40896
rect 0 40838 3299 40840
rect 0 40748 800 40838
rect 3233 40835 3299 40838
rect 68093 40898 68159 40901
rect 69200 40898 70000 40988
rect 68093 40896 70000 40898
rect 68093 40840 68098 40896
rect 68154 40840 70000 40896
rect 68093 40838 70000 40840
rect 68093 40835 68159 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 65648 40832 65968 40833
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 40767 65968 40768
rect 69200 40748 70000 40838
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 50288 40288 50608 40289
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 40223 50608 40224
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 65648 39744 65968 39745
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 39679 65968 39680
rect 0 39538 800 39628
rect 2773 39538 2839 39541
rect 0 39536 2839 39538
rect 0 39480 2778 39536
rect 2834 39480 2839 39536
rect 0 39478 2839 39480
rect 0 39388 800 39478
rect 2773 39475 2839 39478
rect 67265 39538 67331 39541
rect 69200 39538 70000 39628
rect 67265 39536 70000 39538
rect 67265 39480 67270 39536
rect 67326 39480 70000 39536
rect 67265 39478 70000 39480
rect 67265 39475 67331 39478
rect 45645 39402 45711 39405
rect 46749 39402 46815 39405
rect 45645 39400 46815 39402
rect 45645 39344 45650 39400
rect 45706 39344 46754 39400
rect 46810 39344 46815 39400
rect 69200 39388 70000 39478
rect 45645 39342 46815 39344
rect 45645 39339 45711 39342
rect 46749 39339 46815 39342
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 50288 39200 50608 39201
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 39135 50608 39136
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 65648 38656 65968 38657
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 38591 65968 38592
rect 0 38178 800 38268
rect 3233 38178 3299 38181
rect 0 38176 3299 38178
rect 0 38120 3238 38176
rect 3294 38120 3299 38176
rect 0 38118 3299 38120
rect 0 38028 800 38118
rect 3233 38115 3299 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 50288 38112 50608 38113
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 38047 50608 38048
rect 69200 38028 70000 38268
rect 38745 37906 38811 37909
rect 39941 37906 40007 37909
rect 38745 37904 40007 37906
rect 38745 37848 38750 37904
rect 38806 37848 39946 37904
rect 40002 37848 40007 37904
rect 38745 37846 40007 37848
rect 38745 37843 38811 37846
rect 39941 37843 40007 37846
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 65648 37568 65968 37569
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 37503 65968 37504
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 50288 37024 50608 37025
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 36959 50608 36960
rect 0 36818 800 36908
rect 3233 36818 3299 36821
rect 0 36816 3299 36818
rect 0 36760 3238 36816
rect 3294 36760 3299 36816
rect 0 36758 3299 36760
rect 0 36668 800 36758
rect 3233 36755 3299 36758
rect 32305 36682 32371 36685
rect 34881 36682 34947 36685
rect 32305 36680 34947 36682
rect 32305 36624 32310 36680
rect 32366 36624 34886 36680
rect 34942 36624 34947 36680
rect 69200 36668 70000 36908
rect 32305 36622 34947 36624
rect 32305 36619 32371 36622
rect 34881 36619 34947 36622
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 65648 36480 65968 36481
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 36415 65968 36416
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 50288 35936 50608 35937
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 35871 50608 35872
rect 0 35458 800 35548
rect 2773 35458 2839 35461
rect 0 35456 2839 35458
rect 0 35400 2778 35456
rect 2834 35400 2839 35456
rect 0 35398 2839 35400
rect 0 35308 800 35398
rect 2773 35395 2839 35398
rect 67541 35458 67607 35461
rect 69200 35458 70000 35548
rect 67541 35456 70000 35458
rect 67541 35400 67546 35456
rect 67602 35400 70000 35456
rect 67541 35398 70000 35400
rect 67541 35395 67607 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 65648 35392 65968 35393
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 35327 65968 35328
rect 69200 35308 70000 35398
rect 35617 35186 35683 35189
rect 35574 35184 35683 35186
rect 35574 35128 35622 35184
rect 35678 35128 35683 35184
rect 35574 35123 35683 35128
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 35574 34781 35634 35123
rect 50288 34848 50608 34849
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 34783 50608 34784
rect 35574 34776 35683 34781
rect 35574 34720 35622 34776
rect 35678 34720 35683 34776
rect 35574 34718 35683 34720
rect 35617 34715 35683 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 65648 34304 65968 34305
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 34239 65968 34240
rect 0 34098 800 34188
rect 1393 34098 1459 34101
rect 0 34096 1459 34098
rect 0 34040 1398 34096
rect 1454 34040 1459 34096
rect 0 34038 1459 34040
rect 0 33948 800 34038
rect 1393 34035 1459 34038
rect 67265 34098 67331 34101
rect 69200 34098 70000 34188
rect 67265 34096 70000 34098
rect 67265 34040 67270 34096
rect 67326 34040 70000 34096
rect 67265 34038 70000 34040
rect 67265 34035 67331 34038
rect 69200 33948 70000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 50288 33760 50608 33761
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 33695 50608 33696
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 65648 33216 65968 33217
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 33151 65968 33152
rect 0 32588 800 32828
rect 68093 32738 68159 32741
rect 69200 32738 70000 32828
rect 68093 32736 70000 32738
rect 68093 32680 68098 32736
rect 68154 32680 70000 32736
rect 68093 32678 70000 32680
rect 68093 32675 68159 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 50288 32672 50608 32673
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 32607 50608 32608
rect 69200 32588 70000 32678
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 65648 32128 65968 32129
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 32063 65968 32064
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 50288 31584 50608 31585
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 31519 50608 31520
rect 0 31378 800 31468
rect 2773 31378 2839 31381
rect 0 31376 2839 31378
rect 0 31320 2778 31376
rect 2834 31320 2839 31376
rect 0 31318 2839 31320
rect 0 31228 800 31318
rect 2773 31315 2839 31318
rect 67541 31378 67607 31381
rect 69200 31378 70000 31468
rect 67541 31376 70000 31378
rect 67541 31320 67546 31376
rect 67602 31320 70000 31376
rect 67541 31318 70000 31320
rect 67541 31315 67607 31318
rect 69200 31228 70000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 65648 31040 65968 31041
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 30975 65968 30976
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 50288 30496 50608 30497
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 30431 50608 30432
rect 0 30018 800 30108
rect 2865 30018 2931 30021
rect 0 30016 2931 30018
rect 0 29960 2870 30016
rect 2926 29960 2931 30016
rect 0 29958 2931 29960
rect 0 29868 800 29958
rect 2865 29955 2931 29958
rect 66161 30018 66227 30021
rect 69200 30018 70000 30108
rect 66161 30016 70000 30018
rect 66161 29960 66166 30016
rect 66222 29960 70000 30016
rect 66161 29958 70000 29960
rect 66161 29955 66227 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 65648 29952 65968 29953
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 29887 65968 29888
rect 69200 29868 70000 29958
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 50288 29408 50608 29409
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 29343 50608 29344
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 65648 28864 65968 28865
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 28799 65968 28800
rect 0 28508 800 28748
rect 69200 28508 70000 28748
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 50288 28320 50608 28321
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 28255 50608 28256
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 65648 27776 65968 27777
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 27711 65968 27712
rect 0 27298 800 27388
rect 3049 27298 3115 27301
rect 0 27296 3115 27298
rect 0 27240 3054 27296
rect 3110 27240 3115 27296
rect 0 27238 3115 27240
rect 0 27148 800 27238
rect 3049 27235 3115 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 50288 27232 50608 27233
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 27167 50608 27168
rect 69200 27148 70000 27388
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 65648 26688 65968 26689
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 26623 65968 26624
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 50288 26144 50608 26145
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 26079 50608 26080
rect 0 25938 800 26028
rect 2773 25938 2839 25941
rect 0 25936 2839 25938
rect 0 25880 2778 25936
rect 2834 25880 2839 25936
rect 0 25878 2839 25880
rect 0 25788 800 25878
rect 2773 25875 2839 25878
rect 69200 25788 70000 26028
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 65648 25600 65968 25601
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 25535 65968 25536
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 50288 25056 50608 25057
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 24991 50608 24992
rect 0 24578 800 24668
rect 1853 24578 1919 24581
rect 0 24576 1919 24578
rect 0 24520 1858 24576
rect 1914 24520 1919 24576
rect 0 24518 1919 24520
rect 0 24428 800 24518
rect 1853 24515 1919 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 65648 24512 65968 24513
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 24447 65968 24448
rect 69200 24428 70000 24668
rect 0 23898 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 50288 23968 50608 23969
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 23903 50608 23904
rect 2773 23898 2839 23901
rect 0 23896 2839 23898
rect 0 23840 2778 23896
rect 2834 23840 2839 23896
rect 0 23838 2839 23840
rect 0 23748 800 23838
rect 2773 23835 2839 23838
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 65648 23424 65968 23425
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 23359 65968 23360
rect 68093 23218 68159 23221
rect 69200 23218 70000 23308
rect 68093 23216 70000 23218
rect 68093 23160 68098 23216
rect 68154 23160 70000 23216
rect 68093 23158 70000 23160
rect 68093 23155 68159 23158
rect 69200 23068 70000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 50288 22880 50608 22881
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 22815 50608 22816
rect 0 22538 800 22628
rect 2773 22538 2839 22541
rect 0 22536 2839 22538
rect 0 22480 2778 22536
rect 2834 22480 2839 22536
rect 0 22478 2839 22480
rect 0 22388 800 22478
rect 2773 22475 2839 22478
rect 69200 22388 70000 22628
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 65648 22336 65968 22337
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 22271 65968 22272
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 50288 21792 50608 21793
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 21727 50608 21728
rect 0 21178 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 65648 21248 65968 21249
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 21183 65968 21184
rect 1853 21178 1919 21181
rect 0 21176 1919 21178
rect 0 21120 1858 21176
rect 1914 21120 1919 21176
rect 0 21118 1919 21120
rect 0 21028 800 21118
rect 1853 21115 1919 21118
rect 67541 21178 67607 21181
rect 69200 21178 70000 21268
rect 67541 21176 70000 21178
rect 67541 21120 67546 21176
rect 67602 21120 70000 21176
rect 67541 21118 70000 21120
rect 67541 21115 67607 21118
rect 69200 21028 70000 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 50288 20704 50608 20705
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 20639 50608 20640
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 65648 20160 65968 20161
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 20095 65968 20096
rect 0 19668 800 19908
rect 69200 19668 70000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 50288 19616 50608 19617
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 19551 50608 19552
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 65648 19072 65968 19073
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 19007 65968 19008
rect 0 18308 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 50288 18528 50608 18529
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 18463 50608 18464
rect 67817 18458 67883 18461
rect 69200 18458 70000 18548
rect 67817 18456 70000 18458
rect 67817 18400 67822 18456
rect 67878 18400 70000 18456
rect 67817 18398 70000 18400
rect 67817 18395 67883 18398
rect 69200 18308 70000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 65648 17984 65968 17985
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 17919 65968 17920
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 50288 17440 50608 17441
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 17375 50608 17376
rect 0 16948 800 17188
rect 67541 17098 67607 17101
rect 69200 17098 70000 17188
rect 67541 17096 70000 17098
rect 67541 17040 67546 17096
rect 67602 17040 70000 17096
rect 67541 17038 70000 17040
rect 67541 17035 67607 17038
rect 69200 16948 70000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 65648 16896 65968 16897
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 16831 65968 16832
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 50288 16352 50608 16353
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 16287 50608 16288
rect 0 15738 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 65648 15808 65968 15809
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 15743 65968 15744
rect 2957 15738 3023 15741
rect 0 15736 3023 15738
rect 0 15680 2962 15736
rect 3018 15680 3023 15736
rect 0 15678 3023 15680
rect 0 15588 800 15678
rect 2957 15675 3023 15678
rect 66161 15738 66227 15741
rect 69200 15738 70000 15828
rect 66161 15736 70000 15738
rect 66161 15680 66166 15736
rect 66222 15680 70000 15736
rect 66161 15678 70000 15680
rect 66161 15675 66227 15678
rect 69200 15588 70000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 50288 15264 50608 15265
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 15199 50608 15200
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 65648 14720 65968 14721
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 14655 65968 14656
rect 0 14228 800 14468
rect 67541 14378 67607 14381
rect 69200 14378 70000 14468
rect 67541 14376 70000 14378
rect 67541 14320 67546 14376
rect 67602 14320 70000 14376
rect 67541 14318 70000 14320
rect 67541 14315 67607 14318
rect 69200 14228 70000 14318
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 50288 14176 50608 14177
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 14111 50608 14112
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 65648 13632 65968 13633
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 13567 65968 13568
rect 0 13018 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 50288 13088 50608 13089
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 13023 50608 13024
rect 2773 13018 2839 13021
rect 0 13016 2839 13018
rect 0 12960 2778 13016
rect 2834 12960 2839 13016
rect 0 12958 2839 12960
rect 0 12868 800 12958
rect 2773 12955 2839 12958
rect 67817 13018 67883 13021
rect 69200 13018 70000 13108
rect 67817 13016 70000 13018
rect 67817 12960 67822 13016
rect 67878 12960 70000 13016
rect 67817 12958 70000 12960
rect 67817 12955 67883 12958
rect 69200 12868 70000 12958
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 65648 12544 65968 12545
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 12479 65968 12480
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 50288 12000 50608 12001
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 11935 50608 11936
rect 0 11508 800 11748
rect 69200 11508 70000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 65648 11456 65968 11457
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 11391 65968 11392
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 50288 10912 50608 10913
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 10847 50608 10848
rect 0 10148 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 65648 10368 65968 10369
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 10303 65968 10304
rect 69200 10148 70000 10388
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 50288 9824 50608 9825
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 9759 50608 9760
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 65648 9280 65968 9281
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 9215 65968 9216
rect 0 8788 800 9028
rect 69200 8788 70000 9028
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 50288 8736 50608 8737
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 8671 50608 8672
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 65648 8192 65968 8193
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 8127 65968 8128
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 50288 7648 50608 7649
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 7583 50608 7584
rect 1853 7578 1919 7581
rect 0 7576 1919 7578
rect 0 7520 1858 7576
rect 1914 7520 1919 7576
rect 0 7518 1919 7520
rect 0 7428 800 7518
rect 1853 7515 1919 7518
rect 67633 7578 67699 7581
rect 69200 7578 70000 7668
rect 67633 7576 70000 7578
rect 67633 7520 67638 7576
rect 67694 7520 70000 7576
rect 67633 7518 70000 7520
rect 67633 7515 67699 7518
rect 69200 7428 70000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 65648 7104 65968 7105
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 7039 65968 7040
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 50288 6560 50608 6561
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 6495 50608 6496
rect 0 6068 800 6308
rect 67541 6218 67607 6221
rect 69200 6218 70000 6308
rect 67541 6216 70000 6218
rect 67541 6160 67546 6216
rect 67602 6160 70000 6216
rect 67541 6158 70000 6160
rect 67541 6155 67607 6158
rect 69200 6068 70000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 65648 6016 65968 6017
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 5951 65968 5952
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 50288 5472 50608 5473
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 5407 50608 5408
rect 0 4858 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 65648 4928 65968 4929
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 4863 65968 4864
rect 3601 4858 3667 4861
rect 0 4856 3667 4858
rect 0 4800 3606 4856
rect 3662 4800 3667 4856
rect 0 4798 3667 4800
rect 0 4708 800 4798
rect 3601 4795 3667 4798
rect 67541 4858 67607 4861
rect 69200 4858 70000 4948
rect 67541 4856 70000 4858
rect 67541 4800 67546 4856
rect 67602 4800 70000 4856
rect 67541 4798 70000 4800
rect 67541 4795 67607 4798
rect 69200 4708 70000 4798
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 50288 4384 50608 4385
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 4319 50608 4320
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 65648 3840 65968 3841
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 3775 65968 3776
rect 13537 3634 13603 3637
rect 25814 3634 25820 3636
rect 13537 3632 25820 3634
rect 0 3498 800 3588
rect 13537 3576 13542 3632
rect 13598 3576 25820 3632
rect 13537 3574 25820 3576
rect 13537 3571 13603 3574
rect 25814 3572 25820 3574
rect 25884 3572 25890 3636
rect 3141 3498 3207 3501
rect 0 3496 3207 3498
rect 0 3440 3146 3496
rect 3202 3440 3207 3496
rect 0 3438 3207 3440
rect 0 3348 800 3438
rect 3141 3435 3207 3438
rect 4613 3498 4679 3501
rect 25998 3498 26004 3500
rect 4613 3496 26004 3498
rect 4613 3440 4618 3496
rect 4674 3440 26004 3496
rect 4613 3438 26004 3440
rect 4613 3435 4679 3438
rect 25998 3436 26004 3438
rect 26068 3436 26074 3500
rect 69200 3348 70000 3588
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 50288 3296 50608 3297
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 3231 50608 3232
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 65648 2752 65968 2753
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2687 65968 2688
rect 0 2138 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 50288 2208 50608 2209
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2143 50608 2144
rect 2773 2138 2839 2141
rect 0 2136 2839 2138
rect 0 2080 2778 2136
rect 2834 2080 2839 2136
rect 0 2078 2839 2080
rect 0 1988 800 2078
rect 2773 2075 2839 2078
rect 69200 1988 70000 2228
rect 0 778 800 868
rect 2865 778 2931 781
rect 0 776 2931 778
rect 0 720 2870 776
rect 2926 720 2931 776
rect 0 718 2931 720
rect 0 628 800 718
rect 2865 715 2931 718
rect 66161 778 66227 781
rect 69200 778 70000 868
rect 66161 776 70000 778
rect 66161 720 66166 776
rect 66222 720 70000 776
rect 66161 718 70000 720
rect 66161 715 66227 718
rect 69200 628 70000 718
<< via3 >>
rect 19576 69660 19640 69664
rect 19576 69604 19580 69660
rect 19580 69604 19636 69660
rect 19636 69604 19640 69660
rect 19576 69600 19640 69604
rect 19656 69660 19720 69664
rect 19656 69604 19660 69660
rect 19660 69604 19716 69660
rect 19716 69604 19720 69660
rect 19656 69600 19720 69604
rect 19736 69660 19800 69664
rect 19736 69604 19740 69660
rect 19740 69604 19796 69660
rect 19796 69604 19800 69660
rect 19736 69600 19800 69604
rect 19816 69660 19880 69664
rect 19816 69604 19820 69660
rect 19820 69604 19876 69660
rect 19876 69604 19880 69660
rect 19816 69600 19880 69604
rect 50296 69660 50360 69664
rect 50296 69604 50300 69660
rect 50300 69604 50356 69660
rect 50356 69604 50360 69660
rect 50296 69600 50360 69604
rect 50376 69660 50440 69664
rect 50376 69604 50380 69660
rect 50380 69604 50436 69660
rect 50436 69604 50440 69660
rect 50376 69600 50440 69604
rect 50456 69660 50520 69664
rect 50456 69604 50460 69660
rect 50460 69604 50516 69660
rect 50516 69604 50520 69660
rect 50456 69600 50520 69604
rect 50536 69660 50600 69664
rect 50536 69604 50540 69660
rect 50540 69604 50596 69660
rect 50596 69604 50600 69660
rect 50536 69600 50600 69604
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 34936 69116 35000 69120
rect 34936 69060 34940 69116
rect 34940 69060 34996 69116
rect 34996 69060 35000 69116
rect 34936 69056 35000 69060
rect 35016 69116 35080 69120
rect 35016 69060 35020 69116
rect 35020 69060 35076 69116
rect 35076 69060 35080 69116
rect 35016 69056 35080 69060
rect 35096 69116 35160 69120
rect 35096 69060 35100 69116
rect 35100 69060 35156 69116
rect 35156 69060 35160 69116
rect 35096 69056 35160 69060
rect 35176 69116 35240 69120
rect 35176 69060 35180 69116
rect 35180 69060 35236 69116
rect 35236 69060 35240 69116
rect 35176 69056 35240 69060
rect 65656 69116 65720 69120
rect 65656 69060 65660 69116
rect 65660 69060 65716 69116
rect 65716 69060 65720 69116
rect 65656 69056 65720 69060
rect 65736 69116 65800 69120
rect 65736 69060 65740 69116
rect 65740 69060 65796 69116
rect 65796 69060 65800 69116
rect 65736 69056 65800 69060
rect 65816 69116 65880 69120
rect 65816 69060 65820 69116
rect 65820 69060 65876 69116
rect 65876 69060 65880 69116
rect 65816 69056 65880 69060
rect 65896 69116 65960 69120
rect 65896 69060 65900 69116
rect 65900 69060 65956 69116
rect 65956 69060 65960 69116
rect 65896 69056 65960 69060
rect 19576 68572 19640 68576
rect 19576 68516 19580 68572
rect 19580 68516 19636 68572
rect 19636 68516 19640 68572
rect 19576 68512 19640 68516
rect 19656 68572 19720 68576
rect 19656 68516 19660 68572
rect 19660 68516 19716 68572
rect 19716 68516 19720 68572
rect 19656 68512 19720 68516
rect 19736 68572 19800 68576
rect 19736 68516 19740 68572
rect 19740 68516 19796 68572
rect 19796 68516 19800 68572
rect 19736 68512 19800 68516
rect 19816 68572 19880 68576
rect 19816 68516 19820 68572
rect 19820 68516 19876 68572
rect 19876 68516 19880 68572
rect 19816 68512 19880 68516
rect 50296 68572 50360 68576
rect 50296 68516 50300 68572
rect 50300 68516 50356 68572
rect 50356 68516 50360 68572
rect 50296 68512 50360 68516
rect 50376 68572 50440 68576
rect 50376 68516 50380 68572
rect 50380 68516 50436 68572
rect 50436 68516 50440 68572
rect 50376 68512 50440 68516
rect 50456 68572 50520 68576
rect 50456 68516 50460 68572
rect 50460 68516 50516 68572
rect 50516 68516 50520 68572
rect 50456 68512 50520 68516
rect 50536 68572 50600 68576
rect 50536 68516 50540 68572
rect 50540 68516 50596 68572
rect 50596 68516 50600 68572
rect 50536 68512 50600 68516
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 34936 68028 35000 68032
rect 34936 67972 34940 68028
rect 34940 67972 34996 68028
rect 34996 67972 35000 68028
rect 34936 67968 35000 67972
rect 35016 68028 35080 68032
rect 35016 67972 35020 68028
rect 35020 67972 35076 68028
rect 35076 67972 35080 68028
rect 35016 67968 35080 67972
rect 35096 68028 35160 68032
rect 35096 67972 35100 68028
rect 35100 67972 35156 68028
rect 35156 67972 35160 68028
rect 35096 67968 35160 67972
rect 35176 68028 35240 68032
rect 35176 67972 35180 68028
rect 35180 67972 35236 68028
rect 35236 67972 35240 68028
rect 35176 67968 35240 67972
rect 65656 68028 65720 68032
rect 65656 67972 65660 68028
rect 65660 67972 65716 68028
rect 65716 67972 65720 68028
rect 65656 67968 65720 67972
rect 65736 68028 65800 68032
rect 65736 67972 65740 68028
rect 65740 67972 65796 68028
rect 65796 67972 65800 68028
rect 65736 67968 65800 67972
rect 65816 68028 65880 68032
rect 65816 67972 65820 68028
rect 65820 67972 65876 68028
rect 65876 67972 65880 68028
rect 65816 67968 65880 67972
rect 65896 68028 65960 68032
rect 65896 67972 65900 68028
rect 65900 67972 65956 68028
rect 65956 67972 65960 68028
rect 65896 67968 65960 67972
rect 19576 67484 19640 67488
rect 19576 67428 19580 67484
rect 19580 67428 19636 67484
rect 19636 67428 19640 67484
rect 19576 67424 19640 67428
rect 19656 67484 19720 67488
rect 19656 67428 19660 67484
rect 19660 67428 19716 67484
rect 19716 67428 19720 67484
rect 19656 67424 19720 67428
rect 19736 67484 19800 67488
rect 19736 67428 19740 67484
rect 19740 67428 19796 67484
rect 19796 67428 19800 67484
rect 19736 67424 19800 67428
rect 19816 67484 19880 67488
rect 19816 67428 19820 67484
rect 19820 67428 19876 67484
rect 19876 67428 19880 67484
rect 19816 67424 19880 67428
rect 50296 67484 50360 67488
rect 50296 67428 50300 67484
rect 50300 67428 50356 67484
rect 50356 67428 50360 67484
rect 50296 67424 50360 67428
rect 50376 67484 50440 67488
rect 50376 67428 50380 67484
rect 50380 67428 50436 67484
rect 50436 67428 50440 67484
rect 50376 67424 50440 67428
rect 50456 67484 50520 67488
rect 50456 67428 50460 67484
rect 50460 67428 50516 67484
rect 50516 67428 50520 67484
rect 50456 67424 50520 67428
rect 50536 67484 50600 67488
rect 50536 67428 50540 67484
rect 50540 67428 50596 67484
rect 50596 67428 50600 67484
rect 50536 67424 50600 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 34936 66940 35000 66944
rect 34936 66884 34940 66940
rect 34940 66884 34996 66940
rect 34996 66884 35000 66940
rect 34936 66880 35000 66884
rect 35016 66940 35080 66944
rect 35016 66884 35020 66940
rect 35020 66884 35076 66940
rect 35076 66884 35080 66940
rect 35016 66880 35080 66884
rect 35096 66940 35160 66944
rect 35096 66884 35100 66940
rect 35100 66884 35156 66940
rect 35156 66884 35160 66940
rect 35096 66880 35160 66884
rect 35176 66940 35240 66944
rect 35176 66884 35180 66940
rect 35180 66884 35236 66940
rect 35236 66884 35240 66940
rect 35176 66880 35240 66884
rect 65656 66940 65720 66944
rect 65656 66884 65660 66940
rect 65660 66884 65716 66940
rect 65716 66884 65720 66940
rect 65656 66880 65720 66884
rect 65736 66940 65800 66944
rect 65736 66884 65740 66940
rect 65740 66884 65796 66940
rect 65796 66884 65800 66940
rect 65736 66880 65800 66884
rect 65816 66940 65880 66944
rect 65816 66884 65820 66940
rect 65820 66884 65876 66940
rect 65876 66884 65880 66940
rect 65816 66880 65880 66884
rect 65896 66940 65960 66944
rect 65896 66884 65900 66940
rect 65900 66884 65956 66940
rect 65956 66884 65960 66940
rect 65896 66880 65960 66884
rect 19576 66396 19640 66400
rect 19576 66340 19580 66396
rect 19580 66340 19636 66396
rect 19636 66340 19640 66396
rect 19576 66336 19640 66340
rect 19656 66396 19720 66400
rect 19656 66340 19660 66396
rect 19660 66340 19716 66396
rect 19716 66340 19720 66396
rect 19656 66336 19720 66340
rect 19736 66396 19800 66400
rect 19736 66340 19740 66396
rect 19740 66340 19796 66396
rect 19796 66340 19800 66396
rect 19736 66336 19800 66340
rect 19816 66396 19880 66400
rect 19816 66340 19820 66396
rect 19820 66340 19876 66396
rect 19876 66340 19880 66396
rect 19816 66336 19880 66340
rect 50296 66396 50360 66400
rect 50296 66340 50300 66396
rect 50300 66340 50356 66396
rect 50356 66340 50360 66396
rect 50296 66336 50360 66340
rect 50376 66396 50440 66400
rect 50376 66340 50380 66396
rect 50380 66340 50436 66396
rect 50436 66340 50440 66396
rect 50376 66336 50440 66340
rect 50456 66396 50520 66400
rect 50456 66340 50460 66396
rect 50460 66340 50516 66396
rect 50516 66340 50520 66396
rect 50456 66336 50520 66340
rect 50536 66396 50600 66400
rect 50536 66340 50540 66396
rect 50540 66340 50596 66396
rect 50596 66340 50600 66396
rect 50536 66336 50600 66340
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 34936 65852 35000 65856
rect 34936 65796 34940 65852
rect 34940 65796 34996 65852
rect 34996 65796 35000 65852
rect 34936 65792 35000 65796
rect 35016 65852 35080 65856
rect 35016 65796 35020 65852
rect 35020 65796 35076 65852
rect 35076 65796 35080 65852
rect 35016 65792 35080 65796
rect 35096 65852 35160 65856
rect 35096 65796 35100 65852
rect 35100 65796 35156 65852
rect 35156 65796 35160 65852
rect 35096 65792 35160 65796
rect 35176 65852 35240 65856
rect 35176 65796 35180 65852
rect 35180 65796 35236 65852
rect 35236 65796 35240 65852
rect 35176 65792 35240 65796
rect 65656 65852 65720 65856
rect 65656 65796 65660 65852
rect 65660 65796 65716 65852
rect 65716 65796 65720 65852
rect 65656 65792 65720 65796
rect 65736 65852 65800 65856
rect 65736 65796 65740 65852
rect 65740 65796 65796 65852
rect 65796 65796 65800 65852
rect 65736 65792 65800 65796
rect 65816 65852 65880 65856
rect 65816 65796 65820 65852
rect 65820 65796 65876 65852
rect 65876 65796 65880 65852
rect 65816 65792 65880 65796
rect 65896 65852 65960 65856
rect 65896 65796 65900 65852
rect 65900 65796 65956 65852
rect 65956 65796 65960 65852
rect 65896 65792 65960 65796
rect 19576 65308 19640 65312
rect 19576 65252 19580 65308
rect 19580 65252 19636 65308
rect 19636 65252 19640 65308
rect 19576 65248 19640 65252
rect 19656 65308 19720 65312
rect 19656 65252 19660 65308
rect 19660 65252 19716 65308
rect 19716 65252 19720 65308
rect 19656 65248 19720 65252
rect 19736 65308 19800 65312
rect 19736 65252 19740 65308
rect 19740 65252 19796 65308
rect 19796 65252 19800 65308
rect 19736 65248 19800 65252
rect 19816 65308 19880 65312
rect 19816 65252 19820 65308
rect 19820 65252 19876 65308
rect 19876 65252 19880 65308
rect 19816 65248 19880 65252
rect 50296 65308 50360 65312
rect 50296 65252 50300 65308
rect 50300 65252 50356 65308
rect 50356 65252 50360 65308
rect 50296 65248 50360 65252
rect 50376 65308 50440 65312
rect 50376 65252 50380 65308
rect 50380 65252 50436 65308
rect 50436 65252 50440 65308
rect 50376 65248 50440 65252
rect 50456 65308 50520 65312
rect 50456 65252 50460 65308
rect 50460 65252 50516 65308
rect 50516 65252 50520 65308
rect 50456 65248 50520 65252
rect 50536 65308 50600 65312
rect 50536 65252 50540 65308
rect 50540 65252 50596 65308
rect 50596 65252 50600 65308
rect 50536 65248 50600 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 34936 64764 35000 64768
rect 34936 64708 34940 64764
rect 34940 64708 34996 64764
rect 34996 64708 35000 64764
rect 34936 64704 35000 64708
rect 35016 64764 35080 64768
rect 35016 64708 35020 64764
rect 35020 64708 35076 64764
rect 35076 64708 35080 64764
rect 35016 64704 35080 64708
rect 35096 64764 35160 64768
rect 35096 64708 35100 64764
rect 35100 64708 35156 64764
rect 35156 64708 35160 64764
rect 35096 64704 35160 64708
rect 35176 64764 35240 64768
rect 35176 64708 35180 64764
rect 35180 64708 35236 64764
rect 35236 64708 35240 64764
rect 35176 64704 35240 64708
rect 65656 64764 65720 64768
rect 65656 64708 65660 64764
rect 65660 64708 65716 64764
rect 65716 64708 65720 64764
rect 65656 64704 65720 64708
rect 65736 64764 65800 64768
rect 65736 64708 65740 64764
rect 65740 64708 65796 64764
rect 65796 64708 65800 64764
rect 65736 64704 65800 64708
rect 65816 64764 65880 64768
rect 65816 64708 65820 64764
rect 65820 64708 65876 64764
rect 65876 64708 65880 64764
rect 65816 64704 65880 64708
rect 65896 64764 65960 64768
rect 65896 64708 65900 64764
rect 65900 64708 65956 64764
rect 65956 64708 65960 64764
rect 65896 64704 65960 64708
rect 19576 64220 19640 64224
rect 19576 64164 19580 64220
rect 19580 64164 19636 64220
rect 19636 64164 19640 64220
rect 19576 64160 19640 64164
rect 19656 64220 19720 64224
rect 19656 64164 19660 64220
rect 19660 64164 19716 64220
rect 19716 64164 19720 64220
rect 19656 64160 19720 64164
rect 19736 64220 19800 64224
rect 19736 64164 19740 64220
rect 19740 64164 19796 64220
rect 19796 64164 19800 64220
rect 19736 64160 19800 64164
rect 19816 64220 19880 64224
rect 19816 64164 19820 64220
rect 19820 64164 19876 64220
rect 19876 64164 19880 64220
rect 19816 64160 19880 64164
rect 50296 64220 50360 64224
rect 50296 64164 50300 64220
rect 50300 64164 50356 64220
rect 50356 64164 50360 64220
rect 50296 64160 50360 64164
rect 50376 64220 50440 64224
rect 50376 64164 50380 64220
rect 50380 64164 50436 64220
rect 50436 64164 50440 64220
rect 50376 64160 50440 64164
rect 50456 64220 50520 64224
rect 50456 64164 50460 64220
rect 50460 64164 50516 64220
rect 50516 64164 50520 64220
rect 50456 64160 50520 64164
rect 50536 64220 50600 64224
rect 50536 64164 50540 64220
rect 50540 64164 50596 64220
rect 50596 64164 50600 64220
rect 50536 64160 50600 64164
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 34936 63676 35000 63680
rect 34936 63620 34940 63676
rect 34940 63620 34996 63676
rect 34996 63620 35000 63676
rect 34936 63616 35000 63620
rect 35016 63676 35080 63680
rect 35016 63620 35020 63676
rect 35020 63620 35076 63676
rect 35076 63620 35080 63676
rect 35016 63616 35080 63620
rect 35096 63676 35160 63680
rect 35096 63620 35100 63676
rect 35100 63620 35156 63676
rect 35156 63620 35160 63676
rect 35096 63616 35160 63620
rect 35176 63676 35240 63680
rect 35176 63620 35180 63676
rect 35180 63620 35236 63676
rect 35236 63620 35240 63676
rect 35176 63616 35240 63620
rect 65656 63676 65720 63680
rect 65656 63620 65660 63676
rect 65660 63620 65716 63676
rect 65716 63620 65720 63676
rect 65656 63616 65720 63620
rect 65736 63676 65800 63680
rect 65736 63620 65740 63676
rect 65740 63620 65796 63676
rect 65796 63620 65800 63676
rect 65736 63616 65800 63620
rect 65816 63676 65880 63680
rect 65816 63620 65820 63676
rect 65820 63620 65876 63676
rect 65876 63620 65880 63676
rect 65816 63616 65880 63620
rect 65896 63676 65960 63680
rect 65896 63620 65900 63676
rect 65900 63620 65956 63676
rect 65956 63620 65960 63676
rect 65896 63616 65960 63620
rect 19576 63132 19640 63136
rect 19576 63076 19580 63132
rect 19580 63076 19636 63132
rect 19636 63076 19640 63132
rect 19576 63072 19640 63076
rect 19656 63132 19720 63136
rect 19656 63076 19660 63132
rect 19660 63076 19716 63132
rect 19716 63076 19720 63132
rect 19656 63072 19720 63076
rect 19736 63132 19800 63136
rect 19736 63076 19740 63132
rect 19740 63076 19796 63132
rect 19796 63076 19800 63132
rect 19736 63072 19800 63076
rect 19816 63132 19880 63136
rect 19816 63076 19820 63132
rect 19820 63076 19876 63132
rect 19876 63076 19880 63132
rect 19816 63072 19880 63076
rect 50296 63132 50360 63136
rect 50296 63076 50300 63132
rect 50300 63076 50356 63132
rect 50356 63076 50360 63132
rect 50296 63072 50360 63076
rect 50376 63132 50440 63136
rect 50376 63076 50380 63132
rect 50380 63076 50436 63132
rect 50436 63076 50440 63132
rect 50376 63072 50440 63076
rect 50456 63132 50520 63136
rect 50456 63076 50460 63132
rect 50460 63076 50516 63132
rect 50516 63076 50520 63132
rect 50456 63072 50520 63076
rect 50536 63132 50600 63136
rect 50536 63076 50540 63132
rect 50540 63076 50596 63132
rect 50596 63076 50600 63132
rect 50536 63072 50600 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 34936 62588 35000 62592
rect 34936 62532 34940 62588
rect 34940 62532 34996 62588
rect 34996 62532 35000 62588
rect 34936 62528 35000 62532
rect 35016 62588 35080 62592
rect 35016 62532 35020 62588
rect 35020 62532 35076 62588
rect 35076 62532 35080 62588
rect 35016 62528 35080 62532
rect 35096 62588 35160 62592
rect 35096 62532 35100 62588
rect 35100 62532 35156 62588
rect 35156 62532 35160 62588
rect 35096 62528 35160 62532
rect 35176 62588 35240 62592
rect 35176 62532 35180 62588
rect 35180 62532 35236 62588
rect 35236 62532 35240 62588
rect 35176 62528 35240 62532
rect 65656 62588 65720 62592
rect 65656 62532 65660 62588
rect 65660 62532 65716 62588
rect 65716 62532 65720 62588
rect 65656 62528 65720 62532
rect 65736 62588 65800 62592
rect 65736 62532 65740 62588
rect 65740 62532 65796 62588
rect 65796 62532 65800 62588
rect 65736 62528 65800 62532
rect 65816 62588 65880 62592
rect 65816 62532 65820 62588
rect 65820 62532 65876 62588
rect 65876 62532 65880 62588
rect 65816 62528 65880 62532
rect 65896 62588 65960 62592
rect 65896 62532 65900 62588
rect 65900 62532 65956 62588
rect 65956 62532 65960 62588
rect 65896 62528 65960 62532
rect 19576 62044 19640 62048
rect 19576 61988 19580 62044
rect 19580 61988 19636 62044
rect 19636 61988 19640 62044
rect 19576 61984 19640 61988
rect 19656 62044 19720 62048
rect 19656 61988 19660 62044
rect 19660 61988 19716 62044
rect 19716 61988 19720 62044
rect 19656 61984 19720 61988
rect 19736 62044 19800 62048
rect 19736 61988 19740 62044
rect 19740 61988 19796 62044
rect 19796 61988 19800 62044
rect 19736 61984 19800 61988
rect 19816 62044 19880 62048
rect 19816 61988 19820 62044
rect 19820 61988 19876 62044
rect 19876 61988 19880 62044
rect 19816 61984 19880 61988
rect 50296 62044 50360 62048
rect 50296 61988 50300 62044
rect 50300 61988 50356 62044
rect 50356 61988 50360 62044
rect 50296 61984 50360 61988
rect 50376 62044 50440 62048
rect 50376 61988 50380 62044
rect 50380 61988 50436 62044
rect 50436 61988 50440 62044
rect 50376 61984 50440 61988
rect 50456 62044 50520 62048
rect 50456 61988 50460 62044
rect 50460 61988 50516 62044
rect 50516 61988 50520 62044
rect 50456 61984 50520 61988
rect 50536 62044 50600 62048
rect 50536 61988 50540 62044
rect 50540 61988 50596 62044
rect 50596 61988 50600 62044
rect 50536 61984 50600 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 34936 61500 35000 61504
rect 34936 61444 34940 61500
rect 34940 61444 34996 61500
rect 34996 61444 35000 61500
rect 34936 61440 35000 61444
rect 35016 61500 35080 61504
rect 35016 61444 35020 61500
rect 35020 61444 35076 61500
rect 35076 61444 35080 61500
rect 35016 61440 35080 61444
rect 35096 61500 35160 61504
rect 35096 61444 35100 61500
rect 35100 61444 35156 61500
rect 35156 61444 35160 61500
rect 35096 61440 35160 61444
rect 35176 61500 35240 61504
rect 35176 61444 35180 61500
rect 35180 61444 35236 61500
rect 35236 61444 35240 61500
rect 35176 61440 35240 61444
rect 65656 61500 65720 61504
rect 65656 61444 65660 61500
rect 65660 61444 65716 61500
rect 65716 61444 65720 61500
rect 65656 61440 65720 61444
rect 65736 61500 65800 61504
rect 65736 61444 65740 61500
rect 65740 61444 65796 61500
rect 65796 61444 65800 61500
rect 65736 61440 65800 61444
rect 65816 61500 65880 61504
rect 65816 61444 65820 61500
rect 65820 61444 65876 61500
rect 65876 61444 65880 61500
rect 65816 61440 65880 61444
rect 65896 61500 65960 61504
rect 65896 61444 65900 61500
rect 65900 61444 65956 61500
rect 65956 61444 65960 61500
rect 65896 61440 65960 61444
rect 19576 60956 19640 60960
rect 19576 60900 19580 60956
rect 19580 60900 19636 60956
rect 19636 60900 19640 60956
rect 19576 60896 19640 60900
rect 19656 60956 19720 60960
rect 19656 60900 19660 60956
rect 19660 60900 19716 60956
rect 19716 60900 19720 60956
rect 19656 60896 19720 60900
rect 19736 60956 19800 60960
rect 19736 60900 19740 60956
rect 19740 60900 19796 60956
rect 19796 60900 19800 60956
rect 19736 60896 19800 60900
rect 19816 60956 19880 60960
rect 19816 60900 19820 60956
rect 19820 60900 19876 60956
rect 19876 60900 19880 60956
rect 19816 60896 19880 60900
rect 50296 60956 50360 60960
rect 50296 60900 50300 60956
rect 50300 60900 50356 60956
rect 50356 60900 50360 60956
rect 50296 60896 50360 60900
rect 50376 60956 50440 60960
rect 50376 60900 50380 60956
rect 50380 60900 50436 60956
rect 50436 60900 50440 60956
rect 50376 60896 50440 60900
rect 50456 60956 50520 60960
rect 50456 60900 50460 60956
rect 50460 60900 50516 60956
rect 50516 60900 50520 60956
rect 50456 60896 50520 60900
rect 50536 60956 50600 60960
rect 50536 60900 50540 60956
rect 50540 60900 50596 60956
rect 50596 60900 50600 60956
rect 50536 60896 50600 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 65656 60412 65720 60416
rect 65656 60356 65660 60412
rect 65660 60356 65716 60412
rect 65716 60356 65720 60412
rect 65656 60352 65720 60356
rect 65736 60412 65800 60416
rect 65736 60356 65740 60412
rect 65740 60356 65796 60412
rect 65796 60356 65800 60412
rect 65736 60352 65800 60356
rect 65816 60412 65880 60416
rect 65816 60356 65820 60412
rect 65820 60356 65876 60412
rect 65876 60356 65880 60412
rect 65816 60352 65880 60356
rect 65896 60412 65960 60416
rect 65896 60356 65900 60412
rect 65900 60356 65956 60412
rect 65956 60356 65960 60412
rect 65896 60352 65960 60356
rect 19576 59868 19640 59872
rect 19576 59812 19580 59868
rect 19580 59812 19636 59868
rect 19636 59812 19640 59868
rect 19576 59808 19640 59812
rect 19656 59868 19720 59872
rect 19656 59812 19660 59868
rect 19660 59812 19716 59868
rect 19716 59812 19720 59868
rect 19656 59808 19720 59812
rect 19736 59868 19800 59872
rect 19736 59812 19740 59868
rect 19740 59812 19796 59868
rect 19796 59812 19800 59868
rect 19736 59808 19800 59812
rect 19816 59868 19880 59872
rect 19816 59812 19820 59868
rect 19820 59812 19876 59868
rect 19876 59812 19880 59868
rect 19816 59808 19880 59812
rect 50296 59868 50360 59872
rect 50296 59812 50300 59868
rect 50300 59812 50356 59868
rect 50356 59812 50360 59868
rect 50296 59808 50360 59812
rect 50376 59868 50440 59872
rect 50376 59812 50380 59868
rect 50380 59812 50436 59868
rect 50436 59812 50440 59868
rect 50376 59808 50440 59812
rect 50456 59868 50520 59872
rect 50456 59812 50460 59868
rect 50460 59812 50516 59868
rect 50516 59812 50520 59868
rect 50456 59808 50520 59812
rect 50536 59868 50600 59872
rect 50536 59812 50540 59868
rect 50540 59812 50596 59868
rect 50596 59812 50600 59868
rect 50536 59808 50600 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 34936 59324 35000 59328
rect 34936 59268 34940 59324
rect 34940 59268 34996 59324
rect 34996 59268 35000 59324
rect 34936 59264 35000 59268
rect 35016 59324 35080 59328
rect 35016 59268 35020 59324
rect 35020 59268 35076 59324
rect 35076 59268 35080 59324
rect 35016 59264 35080 59268
rect 35096 59324 35160 59328
rect 35096 59268 35100 59324
rect 35100 59268 35156 59324
rect 35156 59268 35160 59324
rect 35096 59264 35160 59268
rect 35176 59324 35240 59328
rect 35176 59268 35180 59324
rect 35180 59268 35236 59324
rect 35236 59268 35240 59324
rect 35176 59264 35240 59268
rect 65656 59324 65720 59328
rect 65656 59268 65660 59324
rect 65660 59268 65716 59324
rect 65716 59268 65720 59324
rect 65656 59264 65720 59268
rect 65736 59324 65800 59328
rect 65736 59268 65740 59324
rect 65740 59268 65796 59324
rect 65796 59268 65800 59324
rect 65736 59264 65800 59268
rect 65816 59324 65880 59328
rect 65816 59268 65820 59324
rect 65820 59268 65876 59324
rect 65876 59268 65880 59324
rect 65816 59264 65880 59268
rect 65896 59324 65960 59328
rect 65896 59268 65900 59324
rect 65900 59268 65956 59324
rect 65956 59268 65960 59324
rect 65896 59264 65960 59268
rect 19576 58780 19640 58784
rect 19576 58724 19580 58780
rect 19580 58724 19636 58780
rect 19636 58724 19640 58780
rect 19576 58720 19640 58724
rect 19656 58780 19720 58784
rect 19656 58724 19660 58780
rect 19660 58724 19716 58780
rect 19716 58724 19720 58780
rect 19656 58720 19720 58724
rect 19736 58780 19800 58784
rect 19736 58724 19740 58780
rect 19740 58724 19796 58780
rect 19796 58724 19800 58780
rect 19736 58720 19800 58724
rect 19816 58780 19880 58784
rect 19816 58724 19820 58780
rect 19820 58724 19876 58780
rect 19876 58724 19880 58780
rect 19816 58720 19880 58724
rect 50296 58780 50360 58784
rect 50296 58724 50300 58780
rect 50300 58724 50356 58780
rect 50356 58724 50360 58780
rect 50296 58720 50360 58724
rect 50376 58780 50440 58784
rect 50376 58724 50380 58780
rect 50380 58724 50436 58780
rect 50436 58724 50440 58780
rect 50376 58720 50440 58724
rect 50456 58780 50520 58784
rect 50456 58724 50460 58780
rect 50460 58724 50516 58780
rect 50516 58724 50520 58780
rect 50456 58720 50520 58724
rect 50536 58780 50600 58784
rect 50536 58724 50540 58780
rect 50540 58724 50596 58780
rect 50596 58724 50600 58780
rect 50536 58720 50600 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 34936 58236 35000 58240
rect 34936 58180 34940 58236
rect 34940 58180 34996 58236
rect 34996 58180 35000 58236
rect 34936 58176 35000 58180
rect 35016 58236 35080 58240
rect 35016 58180 35020 58236
rect 35020 58180 35076 58236
rect 35076 58180 35080 58236
rect 35016 58176 35080 58180
rect 35096 58236 35160 58240
rect 35096 58180 35100 58236
rect 35100 58180 35156 58236
rect 35156 58180 35160 58236
rect 35096 58176 35160 58180
rect 35176 58236 35240 58240
rect 35176 58180 35180 58236
rect 35180 58180 35236 58236
rect 35236 58180 35240 58236
rect 35176 58176 35240 58180
rect 65656 58236 65720 58240
rect 65656 58180 65660 58236
rect 65660 58180 65716 58236
rect 65716 58180 65720 58236
rect 65656 58176 65720 58180
rect 65736 58236 65800 58240
rect 65736 58180 65740 58236
rect 65740 58180 65796 58236
rect 65796 58180 65800 58236
rect 65736 58176 65800 58180
rect 65816 58236 65880 58240
rect 65816 58180 65820 58236
rect 65820 58180 65876 58236
rect 65876 58180 65880 58236
rect 65816 58176 65880 58180
rect 65896 58236 65960 58240
rect 65896 58180 65900 58236
rect 65900 58180 65956 58236
rect 65956 58180 65960 58236
rect 65896 58176 65960 58180
rect 26004 57972 26068 58036
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 65656 57148 65720 57152
rect 65656 57092 65660 57148
rect 65660 57092 65716 57148
rect 65716 57092 65720 57148
rect 65656 57088 65720 57092
rect 65736 57148 65800 57152
rect 65736 57092 65740 57148
rect 65740 57092 65796 57148
rect 65796 57092 65800 57148
rect 65736 57088 65800 57092
rect 65816 57148 65880 57152
rect 65816 57092 65820 57148
rect 65820 57092 65876 57148
rect 65876 57092 65880 57148
rect 65816 57088 65880 57092
rect 65896 57148 65960 57152
rect 65896 57092 65900 57148
rect 65900 57092 65956 57148
rect 65956 57092 65960 57148
rect 65896 57088 65960 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 65656 56060 65720 56064
rect 65656 56004 65660 56060
rect 65660 56004 65716 56060
rect 65716 56004 65720 56060
rect 65656 56000 65720 56004
rect 65736 56060 65800 56064
rect 65736 56004 65740 56060
rect 65740 56004 65796 56060
rect 65796 56004 65800 56060
rect 65736 56000 65800 56004
rect 65816 56060 65880 56064
rect 65816 56004 65820 56060
rect 65820 56004 65876 56060
rect 65876 56004 65880 56060
rect 65816 56000 65880 56004
rect 65896 56060 65960 56064
rect 65896 56004 65900 56060
rect 65900 56004 65956 56060
rect 65956 56004 65960 56060
rect 65896 56000 65960 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 65656 54972 65720 54976
rect 65656 54916 65660 54972
rect 65660 54916 65716 54972
rect 65716 54916 65720 54972
rect 65656 54912 65720 54916
rect 65736 54972 65800 54976
rect 65736 54916 65740 54972
rect 65740 54916 65796 54972
rect 65796 54916 65800 54972
rect 65736 54912 65800 54916
rect 65816 54972 65880 54976
rect 65816 54916 65820 54972
rect 65820 54916 65876 54972
rect 65876 54916 65880 54972
rect 65816 54912 65880 54916
rect 65896 54972 65960 54976
rect 65896 54916 65900 54972
rect 65900 54916 65956 54972
rect 65956 54916 65960 54972
rect 65896 54912 65960 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 65656 53884 65720 53888
rect 65656 53828 65660 53884
rect 65660 53828 65716 53884
rect 65716 53828 65720 53884
rect 65656 53824 65720 53828
rect 65736 53884 65800 53888
rect 65736 53828 65740 53884
rect 65740 53828 65796 53884
rect 65796 53828 65800 53884
rect 65736 53824 65800 53828
rect 65816 53884 65880 53888
rect 65816 53828 65820 53884
rect 65820 53828 65876 53884
rect 65876 53828 65880 53884
rect 65816 53824 65880 53828
rect 65896 53884 65960 53888
rect 65896 53828 65900 53884
rect 65900 53828 65956 53884
rect 65956 53828 65960 53884
rect 65896 53824 65960 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 65656 52796 65720 52800
rect 65656 52740 65660 52796
rect 65660 52740 65716 52796
rect 65716 52740 65720 52796
rect 65656 52736 65720 52740
rect 65736 52796 65800 52800
rect 65736 52740 65740 52796
rect 65740 52740 65796 52796
rect 65796 52740 65800 52796
rect 65736 52736 65800 52740
rect 65816 52796 65880 52800
rect 65816 52740 65820 52796
rect 65820 52740 65876 52796
rect 65876 52740 65880 52796
rect 65816 52736 65880 52740
rect 65896 52796 65960 52800
rect 65896 52740 65900 52796
rect 65900 52740 65956 52796
rect 65956 52740 65960 52796
rect 65896 52736 65960 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 65656 51708 65720 51712
rect 65656 51652 65660 51708
rect 65660 51652 65716 51708
rect 65716 51652 65720 51708
rect 65656 51648 65720 51652
rect 65736 51708 65800 51712
rect 65736 51652 65740 51708
rect 65740 51652 65796 51708
rect 65796 51652 65800 51708
rect 65736 51648 65800 51652
rect 65816 51708 65880 51712
rect 65816 51652 65820 51708
rect 65820 51652 65876 51708
rect 65876 51652 65880 51708
rect 65816 51648 65880 51652
rect 65896 51708 65960 51712
rect 65896 51652 65900 51708
rect 65900 51652 65956 51708
rect 65956 51652 65960 51708
rect 65896 51648 65960 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 65656 50620 65720 50624
rect 65656 50564 65660 50620
rect 65660 50564 65716 50620
rect 65716 50564 65720 50620
rect 65656 50560 65720 50564
rect 65736 50620 65800 50624
rect 65736 50564 65740 50620
rect 65740 50564 65796 50620
rect 65796 50564 65800 50620
rect 65736 50560 65800 50564
rect 65816 50620 65880 50624
rect 65816 50564 65820 50620
rect 65820 50564 65876 50620
rect 65876 50564 65880 50620
rect 65816 50560 65880 50564
rect 65896 50620 65960 50624
rect 65896 50564 65900 50620
rect 65900 50564 65956 50620
rect 65956 50564 65960 50620
rect 65896 50560 65960 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 25820 49736 25884 49740
rect 25820 49680 25870 49736
rect 25870 49680 25884 49736
rect 25820 49676 25884 49680
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 65656 49532 65720 49536
rect 65656 49476 65660 49532
rect 65660 49476 65716 49532
rect 65716 49476 65720 49532
rect 65656 49472 65720 49476
rect 65736 49532 65800 49536
rect 65736 49476 65740 49532
rect 65740 49476 65796 49532
rect 65796 49476 65800 49532
rect 65736 49472 65800 49476
rect 65816 49532 65880 49536
rect 65816 49476 65820 49532
rect 65820 49476 65876 49532
rect 65876 49476 65880 49532
rect 65816 49472 65880 49476
rect 65896 49532 65960 49536
rect 65896 49476 65900 49532
rect 65900 49476 65956 49532
rect 65956 49476 65960 49532
rect 65896 49472 65960 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 65656 48444 65720 48448
rect 65656 48388 65660 48444
rect 65660 48388 65716 48444
rect 65716 48388 65720 48444
rect 65656 48384 65720 48388
rect 65736 48444 65800 48448
rect 65736 48388 65740 48444
rect 65740 48388 65796 48444
rect 65796 48388 65800 48444
rect 65736 48384 65800 48388
rect 65816 48444 65880 48448
rect 65816 48388 65820 48444
rect 65820 48388 65876 48444
rect 65876 48388 65880 48444
rect 65816 48384 65880 48388
rect 65896 48444 65960 48448
rect 65896 48388 65900 48444
rect 65900 48388 65956 48444
rect 65956 48388 65960 48444
rect 65896 48384 65960 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 65656 47356 65720 47360
rect 65656 47300 65660 47356
rect 65660 47300 65716 47356
rect 65716 47300 65720 47356
rect 65656 47296 65720 47300
rect 65736 47356 65800 47360
rect 65736 47300 65740 47356
rect 65740 47300 65796 47356
rect 65796 47300 65800 47356
rect 65736 47296 65800 47300
rect 65816 47356 65880 47360
rect 65816 47300 65820 47356
rect 65820 47300 65876 47356
rect 65876 47300 65880 47356
rect 65816 47296 65880 47300
rect 65896 47356 65960 47360
rect 65896 47300 65900 47356
rect 65900 47300 65956 47356
rect 65956 47300 65960 47356
rect 65896 47296 65960 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 65656 46268 65720 46272
rect 65656 46212 65660 46268
rect 65660 46212 65716 46268
rect 65716 46212 65720 46268
rect 65656 46208 65720 46212
rect 65736 46268 65800 46272
rect 65736 46212 65740 46268
rect 65740 46212 65796 46268
rect 65796 46212 65800 46268
rect 65736 46208 65800 46212
rect 65816 46268 65880 46272
rect 65816 46212 65820 46268
rect 65820 46212 65876 46268
rect 65876 46212 65880 46268
rect 65816 46208 65880 46212
rect 65896 46268 65960 46272
rect 65896 46212 65900 46268
rect 65900 46212 65956 46268
rect 65956 46212 65960 46268
rect 65896 46208 65960 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 65656 45180 65720 45184
rect 65656 45124 65660 45180
rect 65660 45124 65716 45180
rect 65716 45124 65720 45180
rect 65656 45120 65720 45124
rect 65736 45180 65800 45184
rect 65736 45124 65740 45180
rect 65740 45124 65796 45180
rect 65796 45124 65800 45180
rect 65736 45120 65800 45124
rect 65816 45180 65880 45184
rect 65816 45124 65820 45180
rect 65820 45124 65876 45180
rect 65876 45124 65880 45180
rect 65816 45120 65880 45124
rect 65896 45180 65960 45184
rect 65896 45124 65900 45180
rect 65900 45124 65956 45180
rect 65956 45124 65960 45180
rect 65896 45120 65960 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 65656 44092 65720 44096
rect 65656 44036 65660 44092
rect 65660 44036 65716 44092
rect 65716 44036 65720 44092
rect 65656 44032 65720 44036
rect 65736 44092 65800 44096
rect 65736 44036 65740 44092
rect 65740 44036 65796 44092
rect 65796 44036 65800 44092
rect 65736 44032 65800 44036
rect 65816 44092 65880 44096
rect 65816 44036 65820 44092
rect 65820 44036 65876 44092
rect 65876 44036 65880 44092
rect 65816 44032 65880 44036
rect 65896 44092 65960 44096
rect 65896 44036 65900 44092
rect 65900 44036 65956 44092
rect 65956 44036 65960 44092
rect 65896 44032 65960 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 65656 43004 65720 43008
rect 65656 42948 65660 43004
rect 65660 42948 65716 43004
rect 65716 42948 65720 43004
rect 65656 42944 65720 42948
rect 65736 43004 65800 43008
rect 65736 42948 65740 43004
rect 65740 42948 65796 43004
rect 65796 42948 65800 43004
rect 65736 42944 65800 42948
rect 65816 43004 65880 43008
rect 65816 42948 65820 43004
rect 65820 42948 65876 43004
rect 65876 42948 65880 43004
rect 65816 42944 65880 42948
rect 65896 43004 65960 43008
rect 65896 42948 65900 43004
rect 65900 42948 65956 43004
rect 65956 42948 65960 43004
rect 65896 42944 65960 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 65656 41916 65720 41920
rect 65656 41860 65660 41916
rect 65660 41860 65716 41916
rect 65716 41860 65720 41916
rect 65656 41856 65720 41860
rect 65736 41916 65800 41920
rect 65736 41860 65740 41916
rect 65740 41860 65796 41916
rect 65796 41860 65800 41916
rect 65736 41856 65800 41860
rect 65816 41916 65880 41920
rect 65816 41860 65820 41916
rect 65820 41860 65876 41916
rect 65876 41860 65880 41916
rect 65816 41856 65880 41860
rect 65896 41916 65960 41920
rect 65896 41860 65900 41916
rect 65900 41860 65956 41916
rect 65956 41860 65960 41916
rect 65896 41856 65960 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 65656 40828 65720 40832
rect 65656 40772 65660 40828
rect 65660 40772 65716 40828
rect 65716 40772 65720 40828
rect 65656 40768 65720 40772
rect 65736 40828 65800 40832
rect 65736 40772 65740 40828
rect 65740 40772 65796 40828
rect 65796 40772 65800 40828
rect 65736 40768 65800 40772
rect 65816 40828 65880 40832
rect 65816 40772 65820 40828
rect 65820 40772 65876 40828
rect 65876 40772 65880 40828
rect 65816 40768 65880 40772
rect 65896 40828 65960 40832
rect 65896 40772 65900 40828
rect 65900 40772 65956 40828
rect 65956 40772 65960 40828
rect 65896 40768 65960 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 65656 39740 65720 39744
rect 65656 39684 65660 39740
rect 65660 39684 65716 39740
rect 65716 39684 65720 39740
rect 65656 39680 65720 39684
rect 65736 39740 65800 39744
rect 65736 39684 65740 39740
rect 65740 39684 65796 39740
rect 65796 39684 65800 39740
rect 65736 39680 65800 39684
rect 65816 39740 65880 39744
rect 65816 39684 65820 39740
rect 65820 39684 65876 39740
rect 65876 39684 65880 39740
rect 65816 39680 65880 39684
rect 65896 39740 65960 39744
rect 65896 39684 65900 39740
rect 65900 39684 65956 39740
rect 65956 39684 65960 39740
rect 65896 39680 65960 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 65656 38652 65720 38656
rect 65656 38596 65660 38652
rect 65660 38596 65716 38652
rect 65716 38596 65720 38652
rect 65656 38592 65720 38596
rect 65736 38652 65800 38656
rect 65736 38596 65740 38652
rect 65740 38596 65796 38652
rect 65796 38596 65800 38652
rect 65736 38592 65800 38596
rect 65816 38652 65880 38656
rect 65816 38596 65820 38652
rect 65820 38596 65876 38652
rect 65876 38596 65880 38652
rect 65816 38592 65880 38596
rect 65896 38652 65960 38656
rect 65896 38596 65900 38652
rect 65900 38596 65956 38652
rect 65956 38596 65960 38652
rect 65896 38592 65960 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 25820 3572 25884 3636
rect 26004 3436 26068 3500
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 69120 4528 69680
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4528 66944
rect 4208 65856 4528 66880
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 69664 19888 69680
rect 19568 69600 19576 69664
rect 19640 69600 19656 69664
rect 19720 69600 19736 69664
rect 19800 69600 19816 69664
rect 19880 69600 19888 69664
rect 19568 68576 19888 69600
rect 19568 68512 19576 68576
rect 19640 68512 19656 68576
rect 19720 68512 19736 68576
rect 19800 68512 19816 68576
rect 19880 68512 19888 68576
rect 19568 67488 19888 68512
rect 19568 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19888 67488
rect 19568 66400 19888 67424
rect 19568 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19888 66400
rect 19568 65312 19888 66336
rect 19568 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19888 65312
rect 19568 64224 19888 65248
rect 19568 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19888 64224
rect 19568 63136 19888 64160
rect 19568 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19888 63136
rect 19568 62048 19888 63072
rect 19568 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19888 62048
rect 19568 60960 19888 61984
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 59872 19888 60896
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 58784 19888 59808
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 57696 19888 58720
rect 34928 69120 35248 69680
rect 34928 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35248 69120
rect 34928 68032 35248 69056
rect 34928 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35248 68032
rect 34928 66944 35248 67968
rect 34928 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35248 66944
rect 34928 65856 35248 66880
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 64768 35248 65792
rect 34928 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35248 64768
rect 34928 63680 35248 64704
rect 34928 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35248 63680
rect 34928 62592 35248 63616
rect 34928 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35248 62592
rect 34928 61504 35248 62528
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 34928 60416 35248 61440
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 59328 35248 60352
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 58240 35248 59264
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 26003 58036 26069 58037
rect 26003 57972 26004 58036
rect 26068 57972 26069 58036
rect 26003 57971 26069 57972
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 25819 49740 25885 49741
rect 25819 49676 25820 49740
rect 25884 49676 25885 49740
rect 25819 49675 25885 49676
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 25822 3637 25882 49675
rect 25819 3636 25885 3637
rect 25819 3572 25820 3636
rect 25884 3572 25885 3636
rect 25819 3571 25885 3572
rect 26006 3501 26066 57971
rect 34928 57152 35248 58176
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 26003 3500 26069 3501
rect 26003 3436 26004 3500
rect 26068 3436 26069 3500
rect 26003 3435 26069 3436
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 69664 50608 69680
rect 50288 69600 50296 69664
rect 50360 69600 50376 69664
rect 50440 69600 50456 69664
rect 50520 69600 50536 69664
rect 50600 69600 50608 69664
rect 50288 68576 50608 69600
rect 50288 68512 50296 68576
rect 50360 68512 50376 68576
rect 50440 68512 50456 68576
rect 50520 68512 50536 68576
rect 50600 68512 50608 68576
rect 50288 67488 50608 68512
rect 50288 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50608 67488
rect 50288 66400 50608 67424
rect 50288 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50608 66400
rect 50288 65312 50608 66336
rect 50288 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50608 65312
rect 50288 64224 50608 65248
rect 50288 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50608 64224
rect 50288 63136 50608 64160
rect 50288 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50608 63136
rect 50288 62048 50608 63072
rect 50288 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50608 62048
rect 50288 60960 50608 61984
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 59872 50608 60896
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 58784 50608 59808
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 57696 50608 58720
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 69120 65968 69680
rect 65648 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65968 69120
rect 65648 68032 65968 69056
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 66944 65968 67968
rect 65648 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65968 66944
rect 65648 65856 65968 66880
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 64768 65968 65792
rect 65648 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65968 64768
rect 65648 63680 65968 64704
rect 65648 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65968 63680
rect 65648 62592 65968 63616
rect 65648 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65968 62592
rect 65648 61504 65968 62528
rect 65648 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65968 61504
rect 65648 60416 65968 61440
rect 65648 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65968 60416
rect 65648 59328 65968 60352
rect 65648 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65968 59328
rect 65648 58240 65968 59264
rect 65648 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65968 58240
rect 65648 57152 65968 58176
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 56064 65968 57088
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 54976 65968 56000
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 53888 65968 54912
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 52800 65968 53824
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 51712 65968 52736
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 50624 65968 51648
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 49536 65968 50560
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 48448 65968 49472
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 47360 65968 48384
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 46272 65968 47296
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 45184 65968 46208
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 44096 65968 45120
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 43008 65968 44032
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 41920 65968 42944
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 40832 65968 41856
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 39744 65968 40768
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 38656 65968 39680
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 37568 65968 38592
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 28888 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 29808 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 10120 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform -1 0 33304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 20332 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform -1 0 38364 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 20148 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 16928 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1644511149
transform -1 0 67436 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1644511149
transform -1 0 25944 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1644511149
transform -1 0 27048 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1644511149
transform 1 0 25484 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25
timestamp 1644511149
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_33 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1644511149
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_182
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_202
timestamp 1644511149
transform 1 0 19688 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_214
timestamp 1644511149
transform 1 0 20792 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1644511149
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_229
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_236
timestamp 1644511149
transform 1 0 22816 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_342
timestamp 1644511149
transform 1 0 32568 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_354
timestamp 1644511149
transform 1 0 33672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1644511149
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_368
timestamp 1644511149
transform 1 0 34960 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_380
timestamp 1644511149
transform 1 0 36064 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_405
timestamp 1644511149
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1644511149
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1644511149
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_459
timestamp 1644511149
transform 1 0 43332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1644511149
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1644511149
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_489
timestamp 1644511149
transform 1 0 46092 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_493
timestamp 1644511149
transform 1 0 46460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1644511149
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_517
timestamp 1644511149
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1644511149
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_533
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_545
timestamp 1644511149
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1644511149
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_561
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_573
timestamp 1644511149
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1644511149
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_589
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_597
timestamp 1644511149
transform 1 0 56028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_604
timestamp 1644511149
transform 1 0 56672 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_617
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_629
timestamp 1644511149
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1644511149
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_645
timestamp 1644511149
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_657
timestamp 1644511149
transform 1 0 61548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_664
timestamp 1644511149
transform 1 0 62192 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_673
timestamp 1644511149
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_685
timestamp 1644511149
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1644511149
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_707
timestamp 1644511149
transform 1 0 66148 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_715
timestamp 1644511149
transform 1 0 66884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_724
timestamp 1644511149
transform 1 0 67712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_729
timestamp 1644511149
transform 1 0 68172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1644511149
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_97
timestamp 1644511149
transform 1 0 10028 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp 1644511149
transform 1 0 10304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_197
timestamp 1644511149
transform 1 0 19228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1644511149
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_247
timestamp 1644511149
transform 1 0 23828 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_259
timestamp 1644511149
transform 1 0 24932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_271
timestamp 1644511149
transform 1 0 26036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_354
timestamp 1644511149
transform 1 0 33672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1644511149
transform 1 0 35972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_401
timestamp 1644511149
transform 1 0 37996 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_423
timestamp 1644511149
transform 1 0 40020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_435
timestamp 1644511149
transform 1 0 41124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1644511149
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_465
timestamp 1644511149
transform 1 0 43884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_469
timestamp 1644511149
transform 1 0 44252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_494
timestamp 1644511149
transform 1 0 46552 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1644511149
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_517
timestamp 1644511149
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_529
timestamp 1644511149
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_541
timestamp 1644511149
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1644511149
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1644511149
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_573
timestamp 1644511149
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_585
timestamp 1644511149
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_597
timestamp 1644511149
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1644511149
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1644511149
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_617
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_629
timestamp 1644511149
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_641
timestamp 1644511149
transform 1 0 60076 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_668
timestamp 1644511149
transform 1 0 62560 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_673
timestamp 1644511149
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_685
timestamp 1644511149
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_697
timestamp 1644511149
transform 1 0 65228 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_724
timestamp 1644511149
transform 1 0 67712 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_729
timestamp 1644511149
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_12
timestamp 1644511149
transform 1 0 2208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_19
timestamp 1644511149
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_35
timestamp 1644511149
transform 1 0 4324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1644511149
transform 1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_64
timestamp 1644511149
transform 1 0 6992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_71
timestamp 1644511149
transform 1 0 7636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_122
timestamp 1644511149
transform 1 0 12328 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_134
timestamp 1644511149
transform 1 0 13432 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1644511149
transform 1 0 19688 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_214
timestamp 1644511149
transform 1 0 20792 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_226
timestamp 1644511149
transform 1 0 21896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_230
timestamp 1644511149
transform 1 0 22264 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_242
timestamp 1644511149
transform 1 0 23368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1644511149
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_406
timestamp 1644511149
transform 1 0 38456 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1644511149
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_457
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_488
timestamp 1644511149
transform 1 0 46000 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_511
timestamp 1644511149
transform 1 0 48116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_523
timestamp 1644511149
transform 1 0 49220 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1644511149
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1644511149
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1644511149
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1644511149
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1644511149
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1644511149
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1644511149
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_613
timestamp 1644511149
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_625
timestamp 1644511149
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1644511149
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1644511149
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_645
timestamp 1644511149
transform 1 0 60444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_651
timestamp 1644511149
transform 1 0 60996 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_659
timestamp 1644511149
transform 1 0 61732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_682
timestamp 1644511149
transform 1 0 63848 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_694
timestamp 1644511149
transform 1 0 64952 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_701
timestamp 1644511149
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_713
timestamp 1644511149
transform 1 0 66700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_717
timestamp 1644511149
transform 1 0 67068 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_724
timestamp 1644511149
transform 1 0 67712 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_732
timestamp 1644511149
transform 1 0 68448 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_9
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_21
timestamp 1644511149
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_33
timestamp 1644511149
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_46
timestamp 1644511149
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1644511149
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_61
timestamp 1644511149
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_65
timestamp 1644511149
transform 1 0 7084 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_77
timestamp 1644511149
transform 1 0 8188 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_89
timestamp 1644511149
transform 1 0 9292 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_101
timestamp 1644511149
transform 1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1644511149
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_429
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_488
timestamp 1644511149
transform 1 0 46000 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1644511149
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_597
timestamp 1644511149
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1644511149
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1644511149
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_629
timestamp 1644511149
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_641
timestamp 1644511149
transform 1 0 60076 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_647
timestamp 1644511149
transform 1 0 60628 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_651
timestamp 1644511149
transform 1 0 60996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_659
timestamp 1644511149
transform 1 0 61732 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_664
timestamp 1644511149
transform 1 0 62192 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_673
timestamp 1644511149
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_685
timestamp 1644511149
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_697
timestamp 1644511149
transform 1 0 65228 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_724
timestamp 1644511149
transform 1 0 67712 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_729
timestamp 1644511149
transform 1 0 68172 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_63
timestamp 1644511149
transform 1 0 6900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_75
timestamp 1644511149
transform 1 0 8004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_501
timestamp 1644511149
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_513
timestamp 1644511149
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1644511149
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1644511149
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_601
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_613
timestamp 1644511149
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_625
timestamp 1644511149
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1644511149
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1644511149
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_645
timestamp 1644511149
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_657
timestamp 1644511149
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_669
timestamp 1644511149
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_681
timestamp 1644511149
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1644511149
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1644511149
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_701
timestamp 1644511149
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_716
timestamp 1644511149
transform 1 0 66976 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_723
timestamp 1644511149
transform 1 0 67620 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_731
timestamp 1644511149
transform 1 0 68356 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_541
timestamp 1644511149
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1644511149
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_597
timestamp 1644511149
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1644511149
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1644511149
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_629
timestamp 1644511149
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_641
timestamp 1644511149
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_653
timestamp 1644511149
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1644511149
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1644511149
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_673
timestamp 1644511149
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_685
timestamp 1644511149
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_697
timestamp 1644511149
transform 1 0 65228 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_724
timestamp 1644511149
transform 1 0 67712 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_729
timestamp 1644511149
transform 1 0 68172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1644511149
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_613
timestamp 1644511149
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_625
timestamp 1644511149
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1644511149
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1644511149
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_645
timestamp 1644511149
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_657
timestamp 1644511149
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_669
timestamp 1644511149
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_681
timestamp 1644511149
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1644511149
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1644511149
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_701
timestamp 1644511149
transform 1 0 65596 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_707
timestamp 1644511149
transform 1 0 66148 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_711
timestamp 1644511149
transform 1 0 66516 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_718
timestamp 1644511149
transform 1 0 67160 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_725
timestamp 1644511149
transform 1 0 67804 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_529
timestamp 1644511149
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_541
timestamp 1644511149
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1644511149
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1644511149
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_597
timestamp 1644511149
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1644511149
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_617
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_629
timestamp 1644511149
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_641
timestamp 1644511149
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_653
timestamp 1644511149
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1644511149
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1644511149
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_673
timestamp 1644511149
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_685
timestamp 1644511149
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_697
timestamp 1644511149
transform 1 0 65228 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_724
timestamp 1644511149
transform 1 0 67712 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_729
timestamp 1644511149
transform 1 0 68172 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1644511149
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1644511149
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_625
timestamp 1644511149
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1644511149
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1644511149
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_645
timestamp 1644511149
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_657
timestamp 1644511149
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_669
timestamp 1644511149
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_681
timestamp 1644511149
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1644511149
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1644511149
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_701
timestamp 1644511149
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_713
timestamp 1644511149
transform 1 0 66700 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_721
timestamp 1644511149
transform 1 0 67436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_727
timestamp 1644511149
transform 1 0 67988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1644511149
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1644511149
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1644511149
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_629
timestamp 1644511149
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_641
timestamp 1644511149
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_653
timestamp 1644511149
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1644511149
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1644511149
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_673
timestamp 1644511149
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_685
timestamp 1644511149
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_697
timestamp 1644511149
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_709
timestamp 1644511149
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1644511149
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1644511149
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_729
timestamp 1644511149
transform 1 0 68172 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_13
timestamp 1644511149
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1644511149
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1644511149
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_569
timestamp 1644511149
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1644511149
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_625
timestamp 1644511149
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1644511149
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1644511149
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_645
timestamp 1644511149
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_657
timestamp 1644511149
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_669
timestamp 1644511149
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_681
timestamp 1644511149
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1644511149
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1644511149
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_701
timestamp 1644511149
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_713
timestamp 1644511149
transform 1 0 66700 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_721
timestamp 1644511149
transform 1 0 67436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_729
timestamp 1644511149
transform 1 0 68172 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_517
timestamp 1644511149
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_529
timestamp 1644511149
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_541
timestamp 1644511149
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1644511149
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1644511149
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1644511149
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_629
timestamp 1644511149
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_641
timestamp 1644511149
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_653
timestamp 1644511149
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1644511149
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1644511149
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_673
timestamp 1644511149
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_685
timestamp 1644511149
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_697
timestamp 1644511149
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_709
timestamp 1644511149
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1644511149
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1644511149
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_729
timestamp 1644511149
transform 1 0 68172 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1644511149
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1644511149
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_557
timestamp 1644511149
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_569
timestamp 1644511149
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_601
timestamp 1644511149
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_613
timestamp 1644511149
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_625
timestamp 1644511149
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1644511149
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1644511149
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_645
timestamp 1644511149
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_657
timestamp 1644511149
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_669
timestamp 1644511149
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_681
timestamp 1644511149
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1644511149
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1644511149
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_701
timestamp 1644511149
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_713
timestamp 1644511149
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_725
timestamp 1644511149
transform 1 0 67804 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_629
timestamp 1644511149
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_641
timestamp 1644511149
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_653
timestamp 1644511149
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1644511149
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1644511149
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_673
timestamp 1644511149
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_685
timestamp 1644511149
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_697
timestamp 1644511149
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_709
timestamp 1644511149
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1644511149
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1644511149
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_729
timestamp 1644511149
transform 1 0 68172 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1644511149
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_613
timestamp 1644511149
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_625
timestamp 1644511149
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1644511149
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1644511149
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_645
timestamp 1644511149
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_657
timestamp 1644511149
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_669
timestamp 1644511149
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_681
timestamp 1644511149
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1644511149
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1644511149
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_701
timestamp 1644511149
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_713
timestamp 1644511149
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_725
timestamp 1644511149
transform 1 0 67804 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_529
timestamp 1644511149
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_541
timestamp 1644511149
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1644511149
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1644511149
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1644511149
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_629
timestamp 1644511149
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_641
timestamp 1644511149
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_653
timestamp 1644511149
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1644511149
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1644511149
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_673
timestamp 1644511149
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_685
timestamp 1644511149
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_697
timestamp 1644511149
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_709
timestamp 1644511149
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1644511149
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1644511149
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_729
timestamp 1644511149
transform 1 0 68172 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_513
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_557
timestamp 1644511149
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_569
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1644511149
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1644511149
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_625
timestamp 1644511149
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1644511149
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1644511149
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_645
timestamp 1644511149
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_657
timestamp 1644511149
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_669
timestamp 1644511149
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_681
timestamp 1644511149
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1644511149
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1644511149
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_701
timestamp 1644511149
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_713
timestamp 1644511149
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_725
timestamp 1644511149
transform 1 0 67804 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_517
timestamp 1644511149
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_529
timestamp 1644511149
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_541
timestamp 1644511149
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1644511149
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_597
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1644511149
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_629
timestamp 1644511149
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_641
timestamp 1644511149
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_653
timestamp 1644511149
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1644511149
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1644511149
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_673
timestamp 1644511149
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_685
timestamp 1644511149
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_697
timestamp 1644511149
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_709
timestamp 1644511149
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1644511149
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1644511149
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_729
timestamp 1644511149
transform 1 0 68172 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1644511149
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_13
timestamp 1644511149
transform 1 0 2300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1644511149
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1644511149
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1644511149
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_601
timestamp 1644511149
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_613
timestamp 1644511149
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_625
timestamp 1644511149
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1644511149
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1644511149
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_645
timestamp 1644511149
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_657
timestamp 1644511149
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_669
timestamp 1644511149
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_681
timestamp 1644511149
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1644511149
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1644511149
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_701
timestamp 1644511149
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_713
timestamp 1644511149
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_725
timestamp 1644511149
transform 1 0 67804 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_26
timestamp 1644511149
transform 1 0 3496 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_38
timestamp 1644511149
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1644511149
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_346
timestamp 1644511149
transform 1 0 32936 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_350
timestamp 1644511149
transform 1 0 33304 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_362
timestamp 1644511149
transform 1 0 34408 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_374
timestamp 1644511149
transform 1 0 35512 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_386
timestamp 1644511149
transform 1 0 36616 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_517
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_529
timestamp 1644511149
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_541
timestamp 1644511149
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1644511149
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_597
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_629
timestamp 1644511149
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_641
timestamp 1644511149
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_653
timestamp 1644511149
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1644511149
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1644511149
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_673
timestamp 1644511149
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_685
timestamp 1644511149
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_697
timestamp 1644511149
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_709
timestamp 1644511149
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1644511149
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1644511149
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_729
timestamp 1644511149
transform 1 0 68172 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_8
timestamp 1644511149
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1644511149
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1644511149
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1644511149
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_625
timestamp 1644511149
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1644511149
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1644511149
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_645
timestamp 1644511149
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_657
timestamp 1644511149
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_669
timestamp 1644511149
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_681
timestamp 1644511149
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1644511149
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1644511149
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_701
timestamp 1644511149
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_713
timestamp 1644511149
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_729
timestamp 1644511149
transform 1 0 68172 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_541
timestamp 1644511149
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1644511149
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1644511149
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_573
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_585
timestamp 1644511149
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_597
timestamp 1644511149
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1644511149
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_629
timestamp 1644511149
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_641
timestamp 1644511149
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_653
timestamp 1644511149
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1644511149
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1644511149
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_673
timestamp 1644511149
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_685
timestamp 1644511149
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_697
timestamp 1644511149
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_709
timestamp 1644511149
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1644511149
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1644511149
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_729
timestamp 1644511149
transform 1 0 68172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1644511149
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1644511149
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_545
timestamp 1644511149
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_557
timestamp 1644511149
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1644511149
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1644511149
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_601
timestamp 1644511149
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_613
timestamp 1644511149
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_625
timestamp 1644511149
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1644511149
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1644511149
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_645
timestamp 1644511149
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_657
timestamp 1644511149
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_669
timestamp 1644511149
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_681
timestamp 1644511149
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1644511149
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1644511149
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_701
timestamp 1644511149
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_713
timestamp 1644511149
transform 1 0 66700 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_721
timestamp 1644511149
transform 1 0 67436 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_727
timestamp 1644511149
transform 1 0 67988 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_517
timestamp 1644511149
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_529
timestamp 1644511149
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_541
timestamp 1644511149
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1644511149
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1644511149
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_573
timestamp 1644511149
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_585
timestamp 1644511149
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_597
timestamp 1644511149
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1644511149
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_629
timestamp 1644511149
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_641
timestamp 1644511149
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_653
timestamp 1644511149
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1644511149
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1644511149
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_673
timestamp 1644511149
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_685
timestamp 1644511149
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_697
timestamp 1644511149
transform 1 0 65228 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_724
timestamp 1644511149
transform 1 0 67712 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_729
timestamp 1644511149
transform 1 0 68172 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_14
timestamp 1644511149
transform 1 0 2392 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1644511149
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1644511149
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1644511149
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1644511149
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_613
timestamp 1644511149
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_625
timestamp 1644511149
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1644511149
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1644511149
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_645
timestamp 1644511149
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_657
timestamp 1644511149
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_669
timestamp 1644511149
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_681
timestamp 1644511149
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1644511149
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1644511149
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_701
timestamp 1644511149
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_713
timestamp 1644511149
transform 1 0 66700 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_721
timestamp 1644511149
transform 1 0 67436 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_725
timestamp 1644511149
transform 1 0 67804 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_31
timestamp 1644511149
transform 1 0 3956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_43
timestamp 1644511149
transform 1 0 5060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_517
timestamp 1644511149
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1644511149
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1644511149
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_629
timestamp 1644511149
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_641
timestamp 1644511149
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_653
timestamp 1644511149
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1644511149
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1644511149
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_673
timestamp 1644511149
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_685
timestamp 1644511149
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_697
timestamp 1644511149
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_709
timestamp 1644511149
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 1644511149
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 1644511149
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_729
timestamp 1644511149
transform 1 0 68172 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_501
timestamp 1644511149
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_513
timestamp 1644511149
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1644511149
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1644511149
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_557
timestamp 1644511149
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_569
timestamp 1644511149
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_625
timestamp 1644511149
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1644511149
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1644511149
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_645
timestamp 1644511149
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_657
timestamp 1644511149
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_669
timestamp 1644511149
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_681
timestamp 1644511149
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1644511149
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1644511149
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_701
timestamp 1644511149
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_713
timestamp 1644511149
transform 1 0 66700 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_721
timestamp 1644511149
transform 1 0 67436 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_725
timestamp 1644511149
transform 1 0 67804 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_529
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1644511149
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1644511149
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1644511149
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_629
timestamp 1644511149
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_641
timestamp 1644511149
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_653
timestamp 1644511149
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1644511149
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1644511149
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_673
timestamp 1644511149
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_685
timestamp 1644511149
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_697
timestamp 1644511149
transform 1 0 65228 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_724
timestamp 1644511149
transform 1 0 67712 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_729
timestamp 1644511149
transform 1 0 68172 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_513
timestamp 1644511149
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1644511149
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1644511149
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_569
timestamp 1644511149
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1644511149
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_613
timestamp 1644511149
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_625
timestamp 1644511149
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1644511149
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1644511149
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_645
timestamp 1644511149
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_657
timestamp 1644511149
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_669
timestamp 1644511149
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_681
timestamp 1644511149
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1644511149
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1644511149
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_701
timestamp 1644511149
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_713
timestamp 1644511149
transform 1 0 66700 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_721
timestamp 1644511149
transform 1 0 67436 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_727
timestamp 1644511149
transform 1 0 67988 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_290
timestamp 1644511149
transform 1 0 27784 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_302
timestamp 1644511149
transform 1 0 28888 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_314
timestamp 1644511149
transform 1 0 29992 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_326
timestamp 1644511149
transform 1 0 31096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1644511149
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_529
timestamp 1644511149
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_541
timestamp 1644511149
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1644511149
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1644511149
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_585
timestamp 1644511149
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_597
timestamp 1644511149
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1644511149
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_617
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_629
timestamp 1644511149
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_641
timestamp 1644511149
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_653
timestamp 1644511149
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1644511149
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1644511149
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_673
timestamp 1644511149
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_685
timestamp 1644511149
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_697
timestamp 1644511149
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_709
timestamp 1644511149
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1644511149
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1644511149
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_729
timestamp 1644511149
transform 1 0 68172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_601
timestamp 1644511149
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_613
timestamp 1644511149
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_625
timestamp 1644511149
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1644511149
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1644511149
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_645
timestamp 1644511149
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_657
timestamp 1644511149
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_669
timestamp 1644511149
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_681
timestamp 1644511149
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1644511149
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1644511149
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_701
timestamp 1644511149
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_713
timestamp 1644511149
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_729
timestamp 1644511149
transform 1 0 68172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_517
timestamp 1644511149
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1644511149
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1644511149
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1644511149
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_629
timestamp 1644511149
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_641
timestamp 1644511149
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_653
timestamp 1644511149
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1644511149
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1644511149
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_673
timestamp 1644511149
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_685
timestamp 1644511149
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_697
timestamp 1644511149
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_709
timestamp 1644511149
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1644511149
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1644511149
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_729
timestamp 1644511149
transform 1 0 68172 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_501
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_513
timestamp 1644511149
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1644511149
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1644511149
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_613
timestamp 1644511149
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_625
timestamp 1644511149
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1644511149
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1644511149
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_645
timestamp 1644511149
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_657
timestamp 1644511149
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_669
timestamp 1644511149
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_681
timestamp 1644511149
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1644511149
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1644511149
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_701
timestamp 1644511149
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_713
timestamp 1644511149
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_725
timestamp 1644511149
transform 1 0 67804 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1644511149
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_629
timestamp 1644511149
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_641
timestamp 1644511149
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_653
timestamp 1644511149
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1644511149
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1644511149
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_673
timestamp 1644511149
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_685
timestamp 1644511149
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_697
timestamp 1644511149
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_709
timestamp 1644511149
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1644511149
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1644511149
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_729
timestamp 1644511149
transform 1 0 68172 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1644511149
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_601
timestamp 1644511149
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_613
timestamp 1644511149
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_625
timestamp 1644511149
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1644511149
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1644511149
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_645
timestamp 1644511149
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_657
timestamp 1644511149
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_669
timestamp 1644511149
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_681
timestamp 1644511149
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1644511149
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1644511149
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_701
timestamp 1644511149
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_713
timestamp 1644511149
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_725
timestamp 1644511149
transform 1 0 67804 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_11
timestamp 1644511149
transform 1 0 2116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_23
timestamp 1644511149
transform 1 0 3220 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_35
timestamp 1644511149
transform 1 0 4324 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_47
timestamp 1644511149
transform 1 0 5428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1644511149
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1644511149
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_617
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_629
timestamp 1644511149
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_641
timestamp 1644511149
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_653
timestamp 1644511149
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1644511149
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1644511149
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_673
timestamp 1644511149
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_685
timestamp 1644511149
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_697
timestamp 1644511149
transform 1 0 65228 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_724
timestamp 1644511149
transform 1 0 67712 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_729
timestamp 1644511149
transform 1 0 68172 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_7
timestamp 1644511149
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_11
timestamp 1644511149
transform 1 0 2116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_18
timestamp 1644511149
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1644511149
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_513
timestamp 1644511149
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1644511149
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1644511149
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_601
timestamp 1644511149
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_613
timestamp 1644511149
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_625
timestamp 1644511149
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1644511149
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1644511149
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_645
timestamp 1644511149
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_657
timestamp 1644511149
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_669
timestamp 1644511149
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_681
timestamp 1644511149
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1644511149
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1644511149
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_701
timestamp 1644511149
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_713
timestamp 1644511149
transform 1 0 66700 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_721
timestamp 1644511149
transform 1 0 67436 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_727
timestamp 1644511149
transform 1 0 67988 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_28
timestamp 1644511149
transform 1 0 3680 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_40
timestamp 1644511149
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1644511149
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_541
timestamp 1644511149
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1644511149
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1644511149
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_561
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_573
timestamp 1644511149
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_585
timestamp 1644511149
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_597
timestamp 1644511149
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1644511149
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1644511149
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_629
timestamp 1644511149
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_641
timestamp 1644511149
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_653
timestamp 1644511149
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1644511149
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1644511149
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_673
timestamp 1644511149
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_685
timestamp 1644511149
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_697
timestamp 1644511149
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_709
timestamp 1644511149
transform 1 0 66332 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_717
timestamp 1644511149
transform 1 0 67068 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1644511149
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1644511149
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_729
timestamp 1644511149
transform 1 0 68172 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1644511149
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1644511149
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_625
timestamp 1644511149
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1644511149
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1644511149
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_645
timestamp 1644511149
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_657
timestamp 1644511149
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_669
timestamp 1644511149
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_681
timestamp 1644511149
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1644511149
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1644511149
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_701
timestamp 1644511149
transform 1 0 65596 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_707
timestamp 1644511149
transform 1 0 66148 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_729
timestamp 1644511149
transform 1 0 68172 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_517
timestamp 1644511149
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_529
timestamp 1644511149
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_541
timestamp 1644511149
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1644511149
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1644511149
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_597
timestamp 1644511149
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_629
timestamp 1644511149
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_641
timestamp 1644511149
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_653
timestamp 1644511149
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1644511149
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1644511149
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_673
timestamp 1644511149
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_685
timestamp 1644511149
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_697
timestamp 1644511149
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_709
timestamp 1644511149
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_724
timestamp 1644511149
transform 1 0 67712 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_729
timestamp 1644511149
transform 1 0 68172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1644511149
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_337
timestamp 1644511149
transform 1 0 32108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_341
timestamp 1644511149
transform 1 0 32476 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_353
timestamp 1644511149
transform 1 0 33580 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1644511149
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_513
timestamp 1644511149
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1644511149
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1644511149
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_601
timestamp 1644511149
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_613
timestamp 1644511149
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_625
timestamp 1644511149
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1644511149
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1644511149
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_645
timestamp 1644511149
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_657
timestamp 1644511149
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_669
timestamp 1644511149
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_681
timestamp 1644511149
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1644511149
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1644511149
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_701
timestamp 1644511149
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_713
timestamp 1644511149
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_725
timestamp 1644511149
transform 1 0 67804 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_11
timestamp 1644511149
transform 1 0 2116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_19
timestamp 1644511149
transform 1 0 2852 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_26
timestamp 1644511149
transform 1 0 3496 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_38
timestamp 1644511149
transform 1 0 4600 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_50
timestamp 1644511149
transform 1 0 5704 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_325
timestamp 1644511149
transform 1 0 31004 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1644511149
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_353
timestamp 1644511149
transform 1 0 33580 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_357
timestamp 1644511149
transform 1 0 33948 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_517
timestamp 1644511149
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_529
timestamp 1644511149
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_541
timestamp 1644511149
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1644511149
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1644511149
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_597
timestamp 1644511149
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_617
timestamp 1644511149
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_629
timestamp 1644511149
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_641
timestamp 1644511149
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_653
timestamp 1644511149
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1644511149
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1644511149
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_673
timestamp 1644511149
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_685
timestamp 1644511149
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_697
timestamp 1644511149
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_709
timestamp 1644511149
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1644511149
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1644511149
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_729
timestamp 1644511149
transform 1 0 68172 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_11
timestamp 1644511149
transform 1 0 2116 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_346
timestamp 1644511149
transform 1 0 32936 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_352
timestamp 1644511149
transform 1 0 33488 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_370
timestamp 1644511149
transform 1 0 35144 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_382
timestamp 1644511149
transform 1 0 36248 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_394
timestamp 1644511149
transform 1 0 37352 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_406
timestamp 1644511149
transform 1 0 38456 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_418
timestamp 1644511149
transform 1 0 39560 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1644511149
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1644511149
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1644511149
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_533
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_545
timestamp 1644511149
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_557
timestamp 1644511149
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_569
timestamp 1644511149
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1644511149
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_601
timestamp 1644511149
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_613
timestamp 1644511149
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_625
timestamp 1644511149
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1644511149
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1644511149
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_645
timestamp 1644511149
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_657
timestamp 1644511149
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_669
timestamp 1644511149
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_681
timestamp 1644511149
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1644511149
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1644511149
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_701
timestamp 1644511149
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_713
timestamp 1644511149
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_725
timestamp 1644511149
transform 1 0 67804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_323
timestamp 1644511149
transform 1 0 30820 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_328
timestamp 1644511149
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_340
timestamp 1644511149
transform 1 0 32384 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_352
timestamp 1644511149
transform 1 0 33488 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_370
timestamp 1644511149
transform 1 0 35144 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_382
timestamp 1644511149
transform 1 0 36248 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1644511149
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_517
timestamp 1644511149
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_529
timestamp 1644511149
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_541
timestamp 1644511149
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1644511149
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1644511149
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1644511149
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1644511149
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_617
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_629
timestamp 1644511149
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_641
timestamp 1644511149
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_653
timestamp 1644511149
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1644511149
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1644511149
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_673
timestamp 1644511149
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_685
timestamp 1644511149
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_697
timestamp 1644511149
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_709
timestamp 1644511149
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1644511149
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1644511149
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_729
timestamp 1644511149
transform 1 0 68172 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_10
timestamp 1644511149
transform 1 0 2024 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_22
timestamp 1644511149
transform 1 0 3128 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_285
timestamp 1644511149
transform 1 0 27324 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_290
timestamp 1644511149
transform 1 0 27784 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_302
timestamp 1644511149
transform 1 0 28888 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_325
timestamp 1644511149
transform 1 0 31004 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_342
timestamp 1644511149
transform 1 0 32568 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_351
timestamp 1644511149
transform 1 0 33396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_369
timestamp 1644511149
transform 1 0 35052 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_376
timestamp 1644511149
transform 1 0 35696 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_388
timestamp 1644511149
transform 1 0 36800 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_400
timestamp 1644511149
transform 1 0 37904 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_412
timestamp 1644511149
transform 1 0 39008 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_428
timestamp 1644511149
transform 1 0 40480 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_436
timestamp 1644511149
transform 1 0 41216 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_458
timestamp 1644511149
transform 1 0 43240 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_470
timestamp 1644511149
transform 1 0 44344 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_533
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_545
timestamp 1644511149
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_557
timestamp 1644511149
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_569
timestamp 1644511149
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1644511149
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1644511149
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_601
timestamp 1644511149
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_613
timestamp 1644511149
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_625
timestamp 1644511149
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1644511149
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1644511149
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_645
timestamp 1644511149
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_657
timestamp 1644511149
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_669
timestamp 1644511149
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_681
timestamp 1644511149
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1644511149
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1644511149
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_701
timestamp 1644511149
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_713
timestamp 1644511149
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_725
timestamp 1644511149
transform 1 0 67804 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_256
timestamp 1644511149
transform 1 0 24656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1644511149
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_285
timestamp 1644511149
transform 1 0 27324 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_290
timestamp 1644511149
transform 1 0 27784 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_298
timestamp 1644511149
transform 1 0 28520 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_315
timestamp 1644511149
transform 1 0 30084 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_327
timestamp 1644511149
transform 1 0 31188 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_345
timestamp 1644511149
transform 1 0 32844 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_353
timestamp 1644511149
transform 1 0 33580 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_360
timestamp 1644511149
transform 1 0 34224 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_380
timestamp 1644511149
transform 1 0 36064 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_396
timestamp 1644511149
transform 1 0 37536 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_408
timestamp 1644511149
transform 1 0 38640 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_420
timestamp 1644511149
transform 1 0 39744 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_444
timestamp 1644511149
transform 1 0 41952 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1644511149
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1644511149
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1644511149
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1644511149
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1644511149
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_617
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_629
timestamp 1644511149
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_641
timestamp 1644511149
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_653
timestamp 1644511149
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1644511149
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1644511149
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_673
timestamp 1644511149
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_685
timestamp 1644511149
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_697
timestamp 1644511149
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_709
timestamp 1644511149
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1644511149
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1644511149
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_729
timestamp 1644511149
transform 1 0 68172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_242
timestamp 1644511149
transform 1 0 23368 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1644511149
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_274
timestamp 1644511149
transform 1 0 26312 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_280
timestamp 1644511149
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_297
timestamp 1644511149
transform 1 0 28428 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_313
timestamp 1644511149
transform 1 0 29900 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_323
timestamp 1644511149
transform 1 0 30820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_330
timestamp 1644511149
transform 1 0 31464 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_342
timestamp 1644511149
transform 1 0 32568 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_359
timestamp 1644511149
transform 1 0 34132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_370
timestamp 1644511149
transform 1 0 35144 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_382
timestamp 1644511149
transform 1 0 36248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_390
timestamp 1644511149
transform 1 0 36984 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_429
timestamp 1644511149
transform 1 0 40572 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_435
timestamp 1644511149
transform 1 0 41124 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_447
timestamp 1644511149
transform 1 0 42228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_459
timestamp 1644511149
transform 1 0 43332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_471
timestamp 1644511149
transform 1 0 44436 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1644511149
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1644511149
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_545
timestamp 1644511149
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_557
timestamp 1644511149
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_569
timestamp 1644511149
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1644511149
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1644511149
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_601
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_613
timestamp 1644511149
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_625
timestamp 1644511149
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1644511149
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1644511149
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_645
timestamp 1644511149
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_657
timestamp 1644511149
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_669
timestamp 1644511149
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_681
timestamp 1644511149
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1644511149
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1644511149
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_701
timestamp 1644511149
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_713
timestamp 1644511149
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_725
timestamp 1644511149
transform 1 0 67804 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_259
timestamp 1644511149
transform 1 0 24932 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_270
timestamp 1644511149
transform 1 0 25944 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1644511149
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_284
timestamp 1644511149
transform 1 0 27232 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_297
timestamp 1644511149
transform 1 0 28428 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_306
timestamp 1644511149
transform 1 0 29256 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_314
timestamp 1644511149
transform 1 0 29992 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_352
timestamp 1644511149
transform 1 0 33488 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_368
timestamp 1644511149
transform 1 0 34960 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_376
timestamp 1644511149
transform 1 0 35696 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1644511149
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_409
timestamp 1644511149
transform 1 0 38732 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_426
timestamp 1644511149
transform 1 0 40296 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_440
timestamp 1644511149
transform 1 0 41584 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_517
timestamp 1644511149
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_529
timestamp 1644511149
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_541
timestamp 1644511149
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1644511149
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1644511149
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_561
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_573
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_585
timestamp 1644511149
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_597
timestamp 1644511149
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1644511149
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1644511149
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_617
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_629
timestamp 1644511149
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_641
timestamp 1644511149
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_653
timestamp 1644511149
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1644511149
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1644511149
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_673
timestamp 1644511149
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_685
timestamp 1644511149
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_697
timestamp 1644511149
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_709
timestamp 1644511149
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 1644511149
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 1644511149
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_729
timestamp 1644511149
transform 1 0 68172 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_259
timestamp 1644511149
transform 1 0 24932 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_268
timestamp 1644511149
transform 1 0 25760 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_276
timestamp 1644511149
transform 1 0 26496 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_288
timestamp 1644511149
transform 1 0 27600 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_300
timestamp 1644511149
transform 1 0 28704 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_315
timestamp 1644511149
transform 1 0 30084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_332
timestamp 1644511149
transform 1 0 31648 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_344
timestamp 1644511149
transform 1 0 32752 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_356
timestamp 1644511149
transform 1 0 33856 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_369
timestamp 1644511149
transform 1 0 35052 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_386
timestamp 1644511149
transform 1 0 36616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_406
timestamp 1644511149
transform 1 0 38456 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_418
timestamp 1644511149
transform 1 0 39560 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_449
timestamp 1644511149
transform 1 0 42412 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1644511149
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1644511149
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_533
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_545
timestamp 1644511149
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_557
timestamp 1644511149
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_569
timestamp 1644511149
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1644511149
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1644511149
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_601
timestamp 1644511149
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_613
timestamp 1644511149
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_625
timestamp 1644511149
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1644511149
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1644511149
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_645
timestamp 1644511149
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_657
timestamp 1644511149
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_669
timestamp 1644511149
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_681
timestamp 1644511149
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1644511149
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1644511149
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_701
timestamp 1644511149
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_713
timestamp 1644511149
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_725
timestamp 1644511149
transform 1 0 67804 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_255
timestamp 1644511149
transform 1 0 24564 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_272
timestamp 1644511149
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_304
timestamp 1644511149
transform 1 0 29072 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_312
timestamp 1644511149
transform 1 0 29808 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_316
timestamp 1644511149
transform 1 0 30176 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_320
timestamp 1644511149
transform 1 0 30544 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_358
timestamp 1644511149
transform 1 0 34040 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_366
timestamp 1644511149
transform 1 0 34776 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_374
timestamp 1644511149
transform 1 0 35512 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_381
timestamp 1644511149
transform 1 0 36156 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_389
timestamp 1644511149
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_399
timestamp 1644511149
transform 1 0 37812 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_408
timestamp 1644511149
transform 1 0 38640 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_420
timestamp 1644511149
transform 1 0 39744 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_428
timestamp 1644511149
transform 1 0 40480 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_432
timestamp 1644511149
transform 1 0 40848 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_444
timestamp 1644511149
transform 1 0 41952 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_488
timestamp 1644511149
transform 1 0 46000 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_500
timestamp 1644511149
transform 1 0 47104 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_517
timestamp 1644511149
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_529
timestamp 1644511149
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_541
timestamp 1644511149
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1644511149
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1644511149
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_561
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_573
timestamp 1644511149
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_585
timestamp 1644511149
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_597
timestamp 1644511149
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1644511149
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1644511149
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_617
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_629
timestamp 1644511149
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_641
timestamp 1644511149
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_653
timestamp 1644511149
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1644511149
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1644511149
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_673
timestamp 1644511149
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_685
timestamp 1644511149
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_697
timestamp 1644511149
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_709
timestamp 1644511149
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1644511149
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1644511149
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_729
timestamp 1644511149
transform 1 0 68172 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_7
timestamp 1644511149
transform 1 0 1748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_11
timestamp 1644511149
transform 1 0 2116 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_20
timestamp 1644511149
transform 1 0 2944 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_241
timestamp 1644511149
transform 1 0 23276 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1644511149
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_258
timestamp 1644511149
transform 1 0 24840 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_273
timestamp 1644511149
transform 1 0 26220 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_296
timestamp 1644511149
transform 1 0 28336 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_327
timestamp 1644511149
transform 1 0 31188 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_336
timestamp 1644511149
transform 1 0 32016 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_348
timestamp 1644511149
transform 1 0 33120 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1644511149
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_371
timestamp 1644511149
transform 1 0 35236 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_375
timestamp 1644511149
transform 1 0 35604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_387
timestamp 1644511149
transform 1 0 36708 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_393
timestamp 1644511149
transform 1 0 37260 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_405
timestamp 1644511149
transform 1 0 38364 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_414
timestamp 1644511149
transform 1 0 39192 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_426
timestamp 1644511149
transform 1 0 40296 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_437
timestamp 1644511149
transform 1 0 41308 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_449
timestamp 1644511149
transform 1 0 42412 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_461
timestamp 1644511149
transform 1 0 43516 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_473
timestamp 1644511149
transform 1 0 44620 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_480
timestamp 1644511149
transform 1 0 45264 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_492
timestamp 1644511149
transform 1 0 46368 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_504
timestamp 1644511149
transform 1 0 47472 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_516
timestamp 1644511149
transform 1 0 48576 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_528
timestamp 1644511149
transform 1 0 49680 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_545
timestamp 1644511149
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_557
timestamp 1644511149
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_569
timestamp 1644511149
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1644511149
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1644511149
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_589
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_601
timestamp 1644511149
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_613
timestamp 1644511149
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_625
timestamp 1644511149
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1644511149
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1644511149
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_645
timestamp 1644511149
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_657
timestamp 1644511149
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_669
timestamp 1644511149
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_681
timestamp 1644511149
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1644511149
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1644511149
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_701
timestamp 1644511149
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_713
timestamp 1644511149
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_725
timestamp 1644511149
transform 1 0 67804 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_7
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_29
timestamp 1644511149
transform 1 0 3772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_41
timestamp 1644511149
transform 1 0 4876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 1644511149
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_230
timestamp 1644511149
transform 1 0 22264 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_239
timestamp 1644511149
transform 1 0 23092 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_259
timestamp 1644511149
transform 1 0 24932 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_271
timestamp 1644511149
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_297
timestamp 1644511149
transform 1 0 28428 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_314
timestamp 1644511149
transform 1 0 29992 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_322
timestamp 1644511149
transform 1 0 30728 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_328
timestamp 1644511149
transform 1 0 31280 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_341
timestamp 1644511149
transform 1 0 32476 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_347
timestamp 1644511149
transform 1 0 33028 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_351
timestamp 1644511149
transform 1 0 33396 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_381
timestamp 1644511149
transform 1 0 36156 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1644511149
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_398
timestamp 1644511149
transform 1 0 37720 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_402
timestamp 1644511149
transform 1 0 38088 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_406
timestamp 1644511149
transform 1 0 38456 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_410
timestamp 1644511149
transform 1 0 38824 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_418
timestamp 1644511149
transform 1 0 39560 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_426
timestamp 1644511149
transform 1 0 40296 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_444
timestamp 1644511149
transform 1 0 41952 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_460
timestamp 1644511149
transform 1 0 43424 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_466
timestamp 1644511149
transform 1 0 43976 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_483
timestamp 1644511149
transform 1 0 45540 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_495
timestamp 1644511149
transform 1 0 46644 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_517
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_529
timestamp 1644511149
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_541
timestamp 1644511149
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1644511149
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1644511149
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_561
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_573
timestamp 1644511149
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_585
timestamp 1644511149
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_597
timestamp 1644511149
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1644511149
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1644511149
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_617
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_629
timestamp 1644511149
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_641
timestamp 1644511149
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_653
timestamp 1644511149
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1644511149
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1644511149
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_673
timestamp 1644511149
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_685
timestamp 1644511149
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_697
timestamp 1644511149
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_709
timestamp 1644511149
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1644511149
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1644511149
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_729
timestamp 1644511149
transform 1 0 68172 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_12
timestamp 1644511149
transform 1 0 2208 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1644511149
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_229
timestamp 1644511149
transform 1 0 22172 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_243
timestamp 1644511149
transform 1 0 23460 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_256
timestamp 1644511149
transform 1 0 24656 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_268
timestamp 1644511149
transform 1 0 25760 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_280
timestamp 1644511149
transform 1 0 26864 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_292
timestamp 1644511149
transform 1 0 27968 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_299
timestamp 1644511149
transform 1 0 28612 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_312
timestamp 1644511149
transform 1 0 29808 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_324
timestamp 1644511149
transform 1 0 30912 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_342
timestamp 1644511149
transform 1 0 32568 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_348
timestamp 1644511149
transform 1 0 33120 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_354
timestamp 1644511149
transform 1 0 33672 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1644511149
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_368
timestamp 1644511149
transform 1 0 34960 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_390
timestamp 1644511149
transform 1 0 36984 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_412
timestamp 1644511149
transform 1 0 39008 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_432
timestamp 1644511149
transform 1 0 40848 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_440
timestamp 1644511149
transform 1 0 41584 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_452
timestamp 1644511149
transform 1 0 42688 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_460
timestamp 1644511149
transform 1 0 43424 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1644511149
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1644511149
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_545
timestamp 1644511149
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_557
timestamp 1644511149
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_569
timestamp 1644511149
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1644511149
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1644511149
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_589
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_601
timestamp 1644511149
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_613
timestamp 1644511149
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_625
timestamp 1644511149
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1644511149
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1644511149
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_645
timestamp 1644511149
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_657
timestamp 1644511149
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_669
timestamp 1644511149
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_681
timestamp 1644511149
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1644511149
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1644511149
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_701
timestamp 1644511149
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_713
timestamp 1644511149
transform 1 0 66700 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_721
timestamp 1644511149
transform 1 0 67436 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_725
timestamp 1644511149
transform 1 0 67804 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_242
timestamp 1644511149
transform 1 0 23368 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_254
timestamp 1644511149
transform 1 0 24472 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1644511149
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_286
timestamp 1644511149
transform 1 0 27416 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_295
timestamp 1644511149
transform 1 0 28244 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_307
timestamp 1644511149
transform 1 0 29348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_319
timestamp 1644511149
transform 1 0 30452 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_327
timestamp 1644511149
transform 1 0 31188 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_344
timestamp 1644511149
transform 1 0 32752 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_364
timestamp 1644511149
transform 1 0 34592 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_377
timestamp 1644511149
transform 1 0 35788 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_400
timestamp 1644511149
transform 1 0 37904 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_408
timestamp 1644511149
transform 1 0 38640 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_415
timestamp 1644511149
transform 1 0 39284 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_422
timestamp 1644511149
transform 1 0 39928 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_434
timestamp 1644511149
transform 1 0 41032 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_440
timestamp 1644511149
transform 1 0 41584 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_444
timestamp 1644511149
transform 1 0 41952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_454
timestamp 1644511149
transform 1 0 42872 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_462
timestamp 1644511149
transform 1 0 43608 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_467
timestamp 1644511149
transform 1 0 44068 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_474
timestamp 1644511149
transform 1 0 44712 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_486
timestamp 1644511149
transform 1 0 45816 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_498
timestamp 1644511149
transform 1 0 46920 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_517
timestamp 1644511149
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_529
timestamp 1644511149
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_541
timestamp 1644511149
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1644511149
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1644511149
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_585
timestamp 1644511149
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_597
timestamp 1644511149
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1644511149
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1644511149
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_617
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_629
timestamp 1644511149
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_641
timestamp 1644511149
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_653
timestamp 1644511149
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1644511149
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1644511149
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_673
timestamp 1644511149
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_685
timestamp 1644511149
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_697
timestamp 1644511149
transform 1 0 65228 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_724
timestamp 1644511149
transform 1 0 67712 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_729
timestamp 1644511149
transform 1 0 68172 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_9
timestamp 1644511149
transform 1 0 1932 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1644511149
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_229
timestamp 1644511149
transform 1 0 22172 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_234
timestamp 1644511149
transform 1 0 22632 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_243
timestamp 1644511149
transform 1 0 23460 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_264
timestamp 1644511149
transform 1 0 25392 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_272
timestamp 1644511149
transform 1 0 26128 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_279
timestamp 1644511149
transform 1 0 26772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_291
timestamp 1644511149
transform 1 0 27876 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_303
timestamp 1644511149
transform 1 0 28980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_314
timestamp 1644511149
transform 1 0 29992 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_336
timestamp 1644511149
transform 1 0 32016 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_344
timestamp 1644511149
transform 1 0 32752 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_348
timestamp 1644511149
transform 1 0 33120 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1644511149
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_394
timestamp 1644511149
transform 1 0 37352 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_406
timestamp 1644511149
transform 1 0 38456 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_415
timestamp 1644511149
transform 1 0 39284 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_426
timestamp 1644511149
transform 1 0 40296 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_434
timestamp 1644511149
transform 1 0 41032 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_453
timestamp 1644511149
transform 1 0 42780 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_464
timestamp 1644511149
transform 1 0 43792 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_513
timestamp 1644511149
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1644511149
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1644511149
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_545
timestamp 1644511149
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_557
timestamp 1644511149
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_569
timestamp 1644511149
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1644511149
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1644511149
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_589
timestamp 1644511149
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_601
timestamp 1644511149
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_613
timestamp 1644511149
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_625
timestamp 1644511149
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1644511149
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1644511149
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_645
timestamp 1644511149
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_657
timestamp 1644511149
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_669
timestamp 1644511149
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_681
timestamp 1644511149
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1644511149
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1644511149
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_701
timestamp 1644511149
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_713
timestamp 1644511149
transform 1 0 66700 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_721
timestamp 1644511149
transform 1 0 67436 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_727
timestamp 1644511149
transform 1 0 67988 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_247
timestamp 1644511149
transform 1 0 23828 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_259
timestamp 1644511149
transform 1 0 24932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_268
timestamp 1644511149
transform 1 0 25760 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1644511149
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_284
timestamp 1644511149
transform 1 0 27232 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_296
timestamp 1644511149
transform 1 0 28336 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_316
timestamp 1644511149
transform 1 0 30176 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_324
timestamp 1644511149
transform 1 0 30912 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_330
timestamp 1644511149
transform 1 0 31464 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_342
timestamp 1644511149
transform 1 0 32568 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_350
timestamp 1644511149
transform 1 0 33304 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_372
timestamp 1644511149
transform 1 0 35328 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_380
timestamp 1644511149
transform 1 0 36064 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_387
timestamp 1644511149
transform 1 0 36708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_398
timestamp 1644511149
transform 1 0 37720 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_409
timestamp 1644511149
transform 1 0 38732 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_431
timestamp 1644511149
transform 1 0 40756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_435
timestamp 1644511149
transform 1 0 41124 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_440
timestamp 1644511149
transform 1 0 41584 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_457
timestamp 1644511149
transform 1 0 43148 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_465
timestamp 1644511149
transform 1 0 43884 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_475
timestamp 1644511149
transform 1 0 44804 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_495
timestamp 1644511149
transform 1 0 46644 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_517
timestamp 1644511149
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_529
timestamp 1644511149
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_541
timestamp 1644511149
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1644511149
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1644511149
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_561
timestamp 1644511149
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_573
timestamp 1644511149
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_585
timestamp 1644511149
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_597
timestamp 1644511149
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1644511149
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1644511149
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_629
timestamp 1644511149
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_641
timestamp 1644511149
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_653
timestamp 1644511149
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1644511149
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1644511149
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_673
timestamp 1644511149
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_685
timestamp 1644511149
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_697
timestamp 1644511149
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_709
timestamp 1644511149
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_724
timestamp 1644511149
transform 1 0 67712 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_729
timestamp 1644511149
transform 1 0 68172 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_239
timestamp 1644511149
transform 1 0 23092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_263
timestamp 1644511149
transform 1 0 25300 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_271
timestamp 1644511149
transform 1 0 26036 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_298
timestamp 1644511149
transform 1 0 28520 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1644511149
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_312
timestamp 1644511149
transform 1 0 29808 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_327
timestamp 1644511149
transform 1 0 31188 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_339
timestamp 1644511149
transform 1 0 32292 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_356
timestamp 1644511149
transform 1 0 33856 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_370
timestamp 1644511149
transform 1 0 35144 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_390
timestamp 1644511149
transform 1 0 36984 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_399
timestamp 1644511149
transform 1 0 37812 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_407
timestamp 1644511149
transform 1 0 38548 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_411
timestamp 1644511149
transform 1 0 38916 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_456
timestamp 1644511149
transform 1 0 43056 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_464
timestamp 1644511149
transform 1 0 43792 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_472
timestamp 1644511149
transform 1 0 44528 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_495
timestamp 1644511149
transform 1 0 46644 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_517
timestamp 1644511149
transform 1 0 48668 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_529
timestamp 1644511149
transform 1 0 49772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_533
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_545
timestamp 1644511149
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_557
timestamp 1644511149
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_569
timestamp 1644511149
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1644511149
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_601
timestamp 1644511149
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_613
timestamp 1644511149
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_625
timestamp 1644511149
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1644511149
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1644511149
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_645
timestamp 1644511149
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_657
timestamp 1644511149
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_669
timestamp 1644511149
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_681
timestamp 1644511149
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1644511149
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1644511149
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_701
timestamp 1644511149
transform 1 0 65596 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_707
timestamp 1644511149
transform 1 0 66148 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_729
timestamp 1644511149
transform 1 0 68172 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_235
timestamp 1644511149
transform 1 0 22724 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_244
timestamp 1644511149
transform 1 0 23552 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_252
timestamp 1644511149
transform 1 0 24288 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_269
timestamp 1644511149
transform 1 0 25852 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_277
timestamp 1644511149
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_306
timestamp 1644511149
transform 1 0 29256 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_314
timestamp 1644511149
transform 1 0 29992 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_318
timestamp 1644511149
transform 1 0 30360 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_322
timestamp 1644511149
transform 1 0 30728 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1644511149
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_345
timestamp 1644511149
transform 1 0 32844 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_351
timestamp 1644511149
transform 1 0 33396 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_363
timestamp 1644511149
transform 1 0 34500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_371
timestamp 1644511149
transform 1 0 35236 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_382
timestamp 1644511149
transform 1 0 36248 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1644511149
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_401
timestamp 1644511149
transform 1 0 37996 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_407
timestamp 1644511149
transform 1 0 38548 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_416
timestamp 1644511149
transform 1 0 39376 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_422
timestamp 1644511149
transform 1 0 39928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_431
timestamp 1644511149
transform 1 0 40756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_443
timestamp 1644511149
transform 1 0 41860 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_458
timestamp 1644511149
transform 1 0 43240 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_478
timestamp 1644511149
transform 1 0 45080 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_490
timestamp 1644511149
transform 1 0 46184 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_496
timestamp 1644511149
transform 1 0 46736 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_500
timestamp 1644511149
transform 1 0 47104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_517
timestamp 1644511149
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_529
timestamp 1644511149
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_541
timestamp 1644511149
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1644511149
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1644511149
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_561
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_573
timestamp 1644511149
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_585
timestamp 1644511149
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_597
timestamp 1644511149
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1644511149
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1644511149
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_617
timestamp 1644511149
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_629
timestamp 1644511149
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_641
timestamp 1644511149
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_653
timestamp 1644511149
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1644511149
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1644511149
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_673
timestamp 1644511149
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_685
timestamp 1644511149
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_697
timestamp 1644511149
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_709
timestamp 1644511149
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_724
timestamp 1644511149
transform 1 0 67712 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_729
timestamp 1644511149
transform 1 0 68172 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_229
timestamp 1644511149
transform 1 0 22172 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1644511149
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_257
timestamp 1644511149
transform 1 0 24748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_264
timestamp 1644511149
transform 1 0 25392 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_276
timestamp 1644511149
transform 1 0 26496 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_288
timestamp 1644511149
transform 1 0 27600 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_300
timestamp 1644511149
transform 1 0 28704 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_313
timestamp 1644511149
transform 1 0 29900 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_325
timestamp 1644511149
transform 1 0 31004 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_331
timestamp 1644511149
transform 1 0 31556 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_343
timestamp 1644511149
transform 1 0 32660 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_355
timestamp 1644511149
transform 1 0 33764 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_373
timestamp 1644511149
transform 1 0 35420 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_380
timestamp 1644511149
transform 1 0 36064 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_388
timestamp 1644511149
transform 1 0 36800 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_395
timestamp 1644511149
transform 1 0 37444 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_415
timestamp 1644511149
transform 1 0 39284 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_443
timestamp 1644511149
transform 1 0 41860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_449
timestamp 1644511149
transform 1 0 42412 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_466
timestamp 1644511149
transform 1 0 43976 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_474
timestamp 1644511149
transform 1 0 44712 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_486
timestamp 1644511149
transform 1 0 45816 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_498
timestamp 1644511149
transform 1 0 46920 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_510
timestamp 1644511149
transform 1 0 48024 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_522
timestamp 1644511149
transform 1 0 49128 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_530
timestamp 1644511149
transform 1 0 49864 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_545
timestamp 1644511149
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_557
timestamp 1644511149
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_569
timestamp 1644511149
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1644511149
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1644511149
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_601
timestamp 1644511149
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_613
timestamp 1644511149
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_625
timestamp 1644511149
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1644511149
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1644511149
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_645
timestamp 1644511149
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_657
timestamp 1644511149
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_669
timestamp 1644511149
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_681
timestamp 1644511149
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1644511149
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1644511149
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_701
timestamp 1644511149
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_713
timestamp 1644511149
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_725
timestamp 1644511149
transform 1 0 67804 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_13
timestamp 1644511149
transform 1 0 2300 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_25
timestamp 1644511149
transform 1 0 3404 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_37
timestamp 1644511149
transform 1 0 4508 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_49
timestamp 1644511149
transform 1 0 5612 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_240
timestamp 1644511149
transform 1 0 23184 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_252
timestamp 1644511149
transform 1 0 24288 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_259
timestamp 1644511149
transform 1 0 24932 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_267
timestamp 1644511149
transform 1 0 25668 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_272
timestamp 1644511149
transform 1 0 26128 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_287
timestamp 1644511149
transform 1 0 27508 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_299
timestamp 1644511149
transform 1 0 28612 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_311
timestamp 1644511149
transform 1 0 29716 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_315
timestamp 1644511149
transform 1 0 30084 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1644511149
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_340
timestamp 1644511149
transform 1 0 32384 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_346
timestamp 1644511149
transform 1 0 32936 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_352
timestamp 1644511149
transform 1 0 33488 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_364
timestamp 1644511149
transform 1 0 34592 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1644511149
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_403
timestamp 1644511149
transform 1 0 38180 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_418
timestamp 1644511149
transform 1 0 39560 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_430
timestamp 1644511149
transform 1 0 40664 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_435
timestamp 1644511149
transform 1 0 41124 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_439
timestamp 1644511149
transform 1 0 41492 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_443
timestamp 1644511149
transform 1 0 41860 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_465
timestamp 1644511149
transform 1 0 43884 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_469
timestamp 1644511149
transform 1 0 44252 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_481
timestamp 1644511149
transform 1 0 45356 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_498
timestamp 1644511149
transform 1 0 46920 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_508
timestamp 1644511149
transform 1 0 47840 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_520
timestamp 1644511149
transform 1 0 48944 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_532
timestamp 1644511149
transform 1 0 50048 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_544
timestamp 1644511149
transform 1 0 51152 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_556
timestamp 1644511149
transform 1 0 52256 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_561
timestamp 1644511149
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_573
timestamp 1644511149
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_585
timestamp 1644511149
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_597
timestamp 1644511149
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1644511149
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1644511149
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_617
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_629
timestamp 1644511149
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_641
timestamp 1644511149
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_653
timestamp 1644511149
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1644511149
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1644511149
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_673
timestamp 1644511149
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_685
timestamp 1644511149
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_697
timestamp 1644511149
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_709
timestamp 1644511149
transform 1 0 66332 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_717
timestamp 1644511149
transform 1 0 67068 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_724
timestamp 1644511149
transform 1 0 67712 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_729
timestamp 1644511149
transform 1 0 68172 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_205
timestamp 1644511149
transform 1 0 19964 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_217
timestamp 1644511149
transform 1 0 21068 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_229
timestamp 1644511149
transform 1 0 22172 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_234
timestamp 1644511149
transform 1 0 22632 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_241
timestamp 1644511149
transform 1 0 23276 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_249
timestamp 1644511149
transform 1 0 24012 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_259
timestamp 1644511149
transform 1 0 24932 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_279
timestamp 1644511149
transform 1 0 26772 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_314
timestamp 1644511149
transform 1 0 29992 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_322
timestamp 1644511149
transform 1 0 30728 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_331
timestamp 1644511149
transform 1 0 31556 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_339
timestamp 1644511149
transform 1 0 32292 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_358
timestamp 1644511149
transform 1 0 34040 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_386
timestamp 1644511149
transform 1 0 36616 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_397
timestamp 1644511149
transform 1 0 37628 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_403
timestamp 1644511149
transform 1 0 38180 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_407
timestamp 1644511149
transform 1 0 38548 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_414
timestamp 1644511149
transform 1 0 39192 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_434
timestamp 1644511149
transform 1 0 41032 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_438
timestamp 1644511149
transform 1 0 41400 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_449
timestamp 1644511149
transform 1 0 42412 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_458
timestamp 1644511149
transform 1 0 43240 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_466
timestamp 1644511149
transform 1 0 43976 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_474
timestamp 1644511149
transform 1 0 44712 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_485
timestamp 1644511149
transform 1 0 45724 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_497
timestamp 1644511149
transform 1 0 46828 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_503
timestamp 1644511149
transform 1 0 47380 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_533
timestamp 1644511149
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_545
timestamp 1644511149
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_557
timestamp 1644511149
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1644511149
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1644511149
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_601
timestamp 1644511149
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_613
timestamp 1644511149
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_625
timestamp 1644511149
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1644511149
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1644511149
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_645
timestamp 1644511149
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_657
timestamp 1644511149
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_669
timestamp 1644511149
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_681
timestamp 1644511149
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1644511149
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1644511149
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_701
timestamp 1644511149
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_713
timestamp 1644511149
transform 1 0 66700 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_724
timestamp 1644511149
transform 1 0 67712 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_732
timestamp 1644511149
transform 1 0 68448 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_12
timestamp 1644511149
transform 1 0 2208 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_24
timestamp 1644511149
transform 1 0 3312 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_36
timestamp 1644511149
transform 1 0 4416 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_48
timestamp 1644511149
transform 1 0 5520 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_203
timestamp 1644511149
transform 1 0 19780 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_207
timestamp 1644511149
transform 1 0 20148 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_211
timestamp 1644511149
transform 1 0 20516 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_219
timestamp 1644511149
transform 1 0 21252 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_242
timestamp 1644511149
transform 1 0 23368 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_250
timestamp 1644511149
transform 1 0 24104 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_267
timestamp 1644511149
transform 1 0 25668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_284
timestamp 1644511149
transform 1 0 27232 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_296
timestamp 1644511149
transform 1 0 28336 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_315
timestamp 1644511149
transform 1 0 30084 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_323
timestamp 1644511149
transform 1 0 30820 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_332
timestamp 1644511149
transform 1 0 31648 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_344
timestamp 1644511149
transform 1 0 32752 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_351
timestamp 1644511149
transform 1 0 33396 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_363
timestamp 1644511149
transform 1 0 34500 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_367
timestamp 1644511149
transform 1 0 34868 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_371
timestamp 1644511149
transform 1 0 35236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_379
timestamp 1644511149
transform 1 0 35972 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_386
timestamp 1644511149
transform 1 0 36616 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_401
timestamp 1644511149
transform 1 0 37996 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_407
timestamp 1644511149
transform 1 0 38548 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_418
timestamp 1644511149
transform 1 0 39560 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_426
timestamp 1644511149
transform 1 0 40296 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_444
timestamp 1644511149
transform 1 0 41952 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_454
timestamp 1644511149
transform 1 0 42872 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_476
timestamp 1644511149
transform 1 0 44896 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_488
timestamp 1644511149
transform 1 0 46000 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_496
timestamp 1644511149
transform 1 0 46736 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_500
timestamp 1644511149
transform 1 0 47104 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_530
timestamp 1644511149
transform 1 0 49864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_542
timestamp 1644511149
transform 1 0 50968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_554
timestamp 1644511149
transform 1 0 52072 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1644511149
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1644511149
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_629
timestamp 1644511149
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_641
timestamp 1644511149
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_653
timestamp 1644511149
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1644511149
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1644511149
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_673
timestamp 1644511149
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_685
timestamp 1644511149
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_697
timestamp 1644511149
transform 1 0 65228 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_724
timestamp 1644511149
transform 1 0 67712 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_729
timestamp 1644511149
transform 1 0 68172 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_229
timestamp 1644511149
transform 1 0 22172 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_246
timestamp 1644511149
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_258
timestamp 1644511149
transform 1 0 24840 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_280
timestamp 1644511149
transform 1 0 26864 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_292
timestamp 1644511149
transform 1 0 27968 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_302
timestamp 1644511149
transform 1 0 28888 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_312
timestamp 1644511149
transform 1 0 29808 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_320
timestamp 1644511149
transform 1 0 30544 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_340
timestamp 1644511149
transform 1 0 32384 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_353
timestamp 1644511149
transform 1 0 33580 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_361
timestamp 1644511149
transform 1 0 34316 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_395
timestamp 1644511149
transform 1 0 37444 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_399
timestamp 1644511149
transform 1 0 37812 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_416
timestamp 1644511149
transform 1 0 39376 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_431
timestamp 1644511149
transform 1 0 40756 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_449
timestamp 1644511149
transform 1 0 42412 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_464
timestamp 1644511149
transform 1 0 43792 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_509
timestamp 1644511149
transform 1 0 47932 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_521
timestamp 1644511149
transform 1 0 49036 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_529
timestamp 1644511149
transform 1 0 49772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1644511149
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1644511149
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1644511149
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1644511149
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_601
timestamp 1644511149
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_613
timestamp 1644511149
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_625
timestamp 1644511149
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1644511149
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1644511149
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_645
timestamp 1644511149
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_657
timestamp 1644511149
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_669
timestamp 1644511149
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_681
timestamp 1644511149
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1644511149
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1644511149
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_701
timestamp 1644511149
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_713
timestamp 1644511149
transform 1 0 66700 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_721
timestamp 1644511149
transform 1 0 67436 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_727
timestamp 1644511149
transform 1 0 67988 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_18
timestamp 1644511149
transform 1 0 2760 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_30
timestamp 1644511149
transform 1 0 3864 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_42
timestamp 1644511149
transform 1 0 4968 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1644511149
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_233
timestamp 1644511149
transform 1 0 22540 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_247
timestamp 1644511149
transform 1 0 23828 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_255
timestamp 1644511149
transform 1 0 24564 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_259
timestamp 1644511149
transform 1 0 24932 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_265
timestamp 1644511149
transform 1 0 25484 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_294
timestamp 1644511149
transform 1 0 28152 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_308
timestamp 1644511149
transform 1 0 29440 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_321
timestamp 1644511149
transform 1 0 30636 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_332
timestamp 1644511149
transform 1 0 31648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_341
timestamp 1644511149
transform 1 0 32476 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_352
timestamp 1644511149
transform 1 0 33488 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_377
timestamp 1644511149
transform 1 0 35788 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_386
timestamp 1644511149
transform 1 0 36616 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_399
timestamp 1644511149
transform 1 0 37812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_408
timestamp 1644511149
transform 1 0 38640 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_433
timestamp 1644511149
transform 1 0 40940 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_444
timestamp 1644511149
transform 1 0 41952 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_453
timestamp 1644511149
transform 1 0 42780 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_470
timestamp 1644511149
transform 1 0 44344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_474
timestamp 1644511149
transform 1 0 44712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_483
timestamp 1644511149
transform 1 0 45540 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_495
timestamp 1644511149
transform 1 0 46644 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_517
timestamp 1644511149
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_529
timestamp 1644511149
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_541
timestamp 1644511149
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1644511149
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1644511149
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_585
timestamp 1644511149
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_597
timestamp 1644511149
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1644511149
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1644511149
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_617
timestamp 1644511149
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_629
timestamp 1644511149
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_641
timestamp 1644511149
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_653
timestamp 1644511149
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1644511149
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1644511149
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_673
timestamp 1644511149
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_685
timestamp 1644511149
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_697
timestamp 1644511149
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_709
timestamp 1644511149
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 1644511149
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 1644511149
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_729
timestamp 1644511149
transform 1 0 68172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1644511149
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_259
timestamp 1644511149
transform 1 0 24932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_279
timestamp 1644511149
transform 1 0 26772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1644511149
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_341
timestamp 1644511149
transform 1 0 32476 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1644511149
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_368
timestamp 1644511149
transform 1 0 34960 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_372
timestamp 1644511149
transform 1 0 35328 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_383
timestamp 1644511149
transform 1 0 36340 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_391
timestamp 1644511149
transform 1 0 37076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_403
timestamp 1644511149
transform 1 0 38180 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_416
timestamp 1644511149
transform 1 0 39376 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_429
timestamp 1644511149
transform 1 0 40572 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_436
timestamp 1644511149
transform 1 0 41216 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_450
timestamp 1644511149
transform 1 0 42504 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_458
timestamp 1644511149
transform 1 0 43240 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_470
timestamp 1644511149
transform 1 0 44344 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_495
timestamp 1644511149
transform 1 0 46644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_504
timestamp 1644511149
transform 1 0 47472 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_516
timestamp 1644511149
transform 1 0 48576 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_528
timestamp 1644511149
transform 1 0 49680 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_533
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_545
timestamp 1644511149
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_557
timestamp 1644511149
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_569
timestamp 1644511149
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1644511149
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1644511149
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_601
timestamp 1644511149
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_613
timestamp 1644511149
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_625
timestamp 1644511149
transform 1 0 58604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_637
timestamp 1644511149
transform 1 0 59708 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_643
timestamp 1644511149
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_645
timestamp 1644511149
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_657
timestamp 1644511149
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_669
timestamp 1644511149
transform 1 0 62652 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_681
timestamp 1644511149
transform 1 0 63756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_693
timestamp 1644511149
transform 1 0 64860 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_699
timestamp 1644511149
transform 1 0 65412 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_701
timestamp 1644511149
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_713
timestamp 1644511149
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_725
timestamp 1644511149
transform 1 0 67804 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_257
timestamp 1644511149
transform 1 0 24748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_265
timestamp 1644511149
transform 1 0 25484 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_288
timestamp 1644511149
transform 1 0 27600 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_300
timestamp 1644511149
transform 1 0 28704 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_306
timestamp 1644511149
transform 1 0 29256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_323
timestamp 1644511149
transform 1 0 30820 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_340
timestamp 1644511149
transform 1 0 32384 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_344
timestamp 1644511149
transform 1 0 32752 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_355
timestamp 1644511149
transform 1 0 33764 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_367
timestamp 1644511149
transform 1 0 34868 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_380
timestamp 1644511149
transform 1 0 36064 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_401
timestamp 1644511149
transform 1 0 37996 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_437
timestamp 1644511149
transform 1 0 41308 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_445
timestamp 1644511149
transform 1 0 42044 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_459
timestamp 1644511149
transform 1 0 43332 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_467
timestamp 1644511149
transform 1 0 44068 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_481
timestamp 1644511149
transform 1 0 45356 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_493
timestamp 1644511149
transform 1 0 46460 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_501
timestamp 1644511149
transform 1 0 47196 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_526
timestamp 1644511149
transform 1 0 49496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_551
timestamp 1644511149
transform 1 0 51796 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1644511149
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_561
timestamp 1644511149
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_573
timestamp 1644511149
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_585
timestamp 1644511149
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_597
timestamp 1644511149
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1644511149
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1644511149
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_617
timestamp 1644511149
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_629
timestamp 1644511149
transform 1 0 58972 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_641
timestamp 1644511149
transform 1 0 60076 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_653
timestamp 1644511149
transform 1 0 61180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_665
timestamp 1644511149
transform 1 0 62284 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_671
timestamp 1644511149
transform 1 0 62836 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_673
timestamp 1644511149
transform 1 0 63020 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_685
timestamp 1644511149
transform 1 0 64124 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_697
timestamp 1644511149
transform 1 0 65228 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_709
timestamp 1644511149
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_721
timestamp 1644511149
transform 1 0 67436 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_727
timestamp 1644511149
transform 1 0 67988 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_729
timestamp 1644511149
transform 1 0 68172 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_66_206
timestamp 1644511149
transform 1 0 20056 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_214
timestamp 1644511149
transform 1 0 20792 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_231
timestamp 1644511149
transform 1 0 22356 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_243
timestamp 1644511149
transform 1 0 23460 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_247
timestamp 1644511149
transform 1 0 23828 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_269
timestamp 1644511149
transform 1 0 25852 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_281
timestamp 1644511149
transform 1 0 26956 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_292
timestamp 1644511149
transform 1 0 27968 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_304
timestamp 1644511149
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_313
timestamp 1644511149
transform 1 0 29900 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_325
timestamp 1644511149
transform 1 0 31004 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_353
timestamp 1644511149
transform 1 0 33580 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_358
timestamp 1644511149
transform 1 0 34040 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_370
timestamp 1644511149
transform 1 0 35144 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_390
timestamp 1644511149
transform 1 0 36984 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_404
timestamp 1644511149
transform 1 0 38272 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_416
timestamp 1644511149
transform 1 0 39376 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_425
timestamp 1644511149
transform 1 0 40204 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_430
timestamp 1644511149
transform 1 0 40664 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_442
timestamp 1644511149
transform 1 0 41768 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_450
timestamp 1644511149
transform 1 0 42504 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_470
timestamp 1644511149
transform 1 0 44344 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_485
timestamp 1644511149
transform 1 0 45724 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_507
timestamp 1644511149
transform 1 0 47748 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_519
timestamp 1644511149
transform 1 0 48852 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1644511149
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_536
timestamp 1644511149
transform 1 0 50416 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_548
timestamp 1644511149
transform 1 0 51520 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_560
timestamp 1644511149
transform 1 0 52624 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_572
timestamp 1644511149
transform 1 0 53728 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_584
timestamp 1644511149
transform 1 0 54832 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_589
timestamp 1644511149
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_601
timestamp 1644511149
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_613
timestamp 1644511149
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_625
timestamp 1644511149
transform 1 0 58604 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_637
timestamp 1644511149
transform 1 0 59708 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_643
timestamp 1644511149
transform 1 0 60260 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_645
timestamp 1644511149
transform 1 0 60444 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_657
timestamp 1644511149
transform 1 0 61548 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_669
timestamp 1644511149
transform 1 0 62652 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_681
timestamp 1644511149
transform 1 0 63756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_693
timestamp 1644511149
transform 1 0 64860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_699
timestamp 1644511149
transform 1 0 65412 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_701
timestamp 1644511149
transform 1 0 65596 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_713
timestamp 1644511149
transform 1 0 66700 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_725
timestamp 1644511149
transform 1 0 67804 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_10
timestamp 1644511149
transform 1 0 2024 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_22
timestamp 1644511149
transform 1 0 3128 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_34
timestamp 1644511149
transform 1 0 4232 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_46
timestamp 1644511149
transform 1 0 5336 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp 1644511149
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_204
timestamp 1644511149
transform 1 0 19872 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_220
timestamp 1644511149
transform 1 0 21344 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_241
timestamp 1644511149
transform 1 0 23276 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_268
timestamp 1644511149
transform 1 0 25760 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1644511149
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_298
timestamp 1644511149
transform 1 0 28520 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_310
timestamp 1644511149
transform 1 0 29624 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_322
timestamp 1644511149
transform 1 0 30728 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_327
timestamp 1644511149
transform 1 0 31188 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_342
timestamp 1644511149
transform 1 0 32568 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_350
timestamp 1644511149
transform 1 0 33304 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_372
timestamp 1644511149
transform 1 0 35328 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_376
timestamp 1644511149
transform 1 0 35696 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_381
timestamp 1644511149
transform 1 0 36156 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_388
timestamp 1644511149
transform 1 0 36800 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_399
timestamp 1644511149
transform 1 0 37812 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_416
timestamp 1644511149
transform 1 0 39376 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_431
timestamp 1644511149
transform 1 0 40756 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_437
timestamp 1644511149
transform 1 0 41308 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_443
timestamp 1644511149
transform 1 0 41860 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_456
timestamp 1644511149
transform 1 0 43056 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_465
timestamp 1644511149
transform 1 0 43884 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_489
timestamp 1644511149
transform 1 0 46092 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_501
timestamp 1644511149
transform 1 0 47196 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_517
timestamp 1644511149
transform 1 0 48668 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_539
timestamp 1644511149
transform 1 0 50692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_551
timestamp 1644511149
transform 1 0 51796 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1644511149
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_561
timestamp 1644511149
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_573
timestamp 1644511149
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_585
timestamp 1644511149
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_597
timestamp 1644511149
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1644511149
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1644511149
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_617
timestamp 1644511149
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_629
timestamp 1644511149
transform 1 0 58972 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_641
timestamp 1644511149
transform 1 0 60076 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_653
timestamp 1644511149
transform 1 0 61180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_665
timestamp 1644511149
transform 1 0 62284 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_671
timestamp 1644511149
transform 1 0 62836 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_673
timestamp 1644511149
transform 1 0 63020 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_685
timestamp 1644511149
transform 1 0 64124 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_697
timestamp 1644511149
transform 1 0 65228 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_709
timestamp 1644511149
transform 1 0 66332 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_721
timestamp 1644511149
transform 1 0 67436 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_727
timestamp 1644511149
transform 1 0 67988 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_729
timestamp 1644511149
transform 1 0 68172 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_24
timestamp 1644511149
transform 1 0 3312 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_219
timestamp 1644511149
transform 1 0 21252 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_231
timestamp 1644511149
transform 1 0 22356 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1644511149
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_261
timestamp 1644511149
transform 1 0 25116 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_270
timestamp 1644511149
transform 1 0 25944 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_278
timestamp 1644511149
transform 1 0 26680 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_286
timestamp 1644511149
transform 1 0 27416 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_292
timestamp 1644511149
transform 1 0 27968 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_298
timestamp 1644511149
transform 1 0 28520 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_306
timestamp 1644511149
transform 1 0 29256 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_315
timestamp 1644511149
transform 1 0 30084 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_322
timestamp 1644511149
transform 1 0 30728 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_344
timestamp 1644511149
transform 1 0 32752 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_356
timestamp 1644511149
transform 1 0 33856 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_369
timestamp 1644511149
transform 1 0 35052 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_375
timestamp 1644511149
transform 1 0 35604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_387
timestamp 1644511149
transform 1 0 36708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_68_398
timestamp 1644511149
transform 1 0 37720 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_68_412
timestamp 1644511149
transform 1 0 39008 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_429
timestamp 1644511149
transform 1 0 40572 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_438
timestamp 1644511149
transform 1 0 41400 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_446
timestamp 1644511149
transform 1 0 42136 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_456
timestamp 1644511149
transform 1 0 43056 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_463
timestamp 1644511149
transform 1 0 43700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_485
timestamp 1644511149
transform 1 0 45724 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_492
timestamp 1644511149
transform 1 0 46368 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_68_521
timestamp 1644511149
transform 1 0 49036 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_529
timestamp 1644511149
transform 1 0 49772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_533
timestamp 1644511149
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_545
timestamp 1644511149
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_557
timestamp 1644511149
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_569
timestamp 1644511149
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1644511149
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1644511149
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_589
timestamp 1644511149
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_601
timestamp 1644511149
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_613
timestamp 1644511149
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_625
timestamp 1644511149
transform 1 0 58604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_637
timestamp 1644511149
transform 1 0 59708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_643
timestamp 1644511149
transform 1 0 60260 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_645
timestamp 1644511149
transform 1 0 60444 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_657
timestamp 1644511149
transform 1 0 61548 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_669
timestamp 1644511149
transform 1 0 62652 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_681
timestamp 1644511149
transform 1 0 63756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_693
timestamp 1644511149
transform 1 0 64860 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_699
timestamp 1644511149
transform 1 0 65412 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_701
timestamp 1644511149
transform 1 0 65596 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_713
timestamp 1644511149
transform 1 0 66700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_725
timestamp 1644511149
transform 1 0 67804 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_7
timestamp 1644511149
transform 1 0 1748 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_19
timestamp 1644511149
transform 1 0 2852 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_31
timestamp 1644511149
transform 1 0 3956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_43
timestamp 1644511149
transform 1 0 5060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_201
timestamp 1644511149
transform 1 0 19596 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1644511149
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_233
timestamp 1644511149
transform 1 0 22540 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_257
timestamp 1644511149
transform 1 0 24748 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_265
timestamp 1644511149
transform 1 0 25484 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_271
timestamp 1644511149
transform 1 0 26036 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_276
timestamp 1644511149
transform 1 0 26496 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_284
timestamp 1644511149
transform 1 0 27232 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_302
timestamp 1644511149
transform 1 0 28888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_322
timestamp 1644511149
transform 1 0 30728 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_328
timestamp 1644511149
transform 1 0 31280 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_332
timestamp 1644511149
transform 1 0 31648 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_342
timestamp 1644511149
transform 1 0 32568 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_348
timestamp 1644511149
transform 1 0 33120 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_370
timestamp 1644511149
transform 1 0 35144 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_382
timestamp 1644511149
transform 1 0 36248 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_390
timestamp 1644511149
transform 1 0 36984 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_398
timestamp 1644511149
transform 1 0 37720 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_406
timestamp 1644511149
transform 1 0 38456 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_410
timestamp 1644511149
transform 1 0 38824 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_415
timestamp 1644511149
transform 1 0 39284 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_421
timestamp 1644511149
transform 1 0 39836 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_438
timestamp 1644511149
transform 1 0 41400 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_446
timestamp 1644511149
transform 1 0 42136 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_455
timestamp 1644511149
transform 1 0 42964 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_463
timestamp 1644511149
transform 1 0 43700 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_480
timestamp 1644511149
transform 1 0 45264 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_488
timestamp 1644511149
transform 1 0 46000 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_505
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_517
timestamp 1644511149
transform 1 0 48668 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_539
timestamp 1644511149
transform 1 0 50692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_551
timestamp 1644511149
transform 1 0 51796 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1644511149
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_561
timestamp 1644511149
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_573
timestamp 1644511149
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_585
timestamp 1644511149
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_597
timestamp 1644511149
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1644511149
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1644511149
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_617
timestamp 1644511149
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_629
timestamp 1644511149
transform 1 0 58972 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_641
timestamp 1644511149
transform 1 0 60076 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_653
timestamp 1644511149
transform 1 0 61180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_665
timestamp 1644511149
transform 1 0 62284 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_671
timestamp 1644511149
transform 1 0 62836 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_673
timestamp 1644511149
transform 1 0 63020 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_685
timestamp 1644511149
transform 1 0 64124 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_697
timestamp 1644511149
transform 1 0 65228 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_709
timestamp 1644511149
transform 1 0 66332 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_717
timestamp 1644511149
transform 1 0 67068 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_724
timestamp 1644511149
transform 1 0 67712 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_729
timestamp 1644511149
transform 1 0 68172 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1644511149
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_192
timestamp 1644511149
transform 1 0 18768 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_218
timestamp 1644511149
transform 1 0 21160 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_230
timestamp 1644511149
transform 1 0 22264 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_238
timestamp 1644511149
transform 1 0 23000 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_244
timestamp 1644511149
transform 1 0 23552 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_269
timestamp 1644511149
transform 1 0 25852 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_298
timestamp 1644511149
transform 1 0 28520 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_306
timestamp 1644511149
transform 1 0 29256 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_313
timestamp 1644511149
transform 1 0 29900 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_325
timestamp 1644511149
transform 1 0 31004 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_337
timestamp 1644511149
transform 1 0 32108 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_349
timestamp 1644511149
transform 1 0 33212 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_361
timestamp 1644511149
transform 1 0 34316 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_369
timestamp 1644511149
transform 1 0 35052 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_375
timestamp 1644511149
transform 1 0 35604 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_381
timestamp 1644511149
transform 1 0 36156 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_385
timestamp 1644511149
transform 1 0 36524 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_395
timestamp 1644511149
transform 1 0 37444 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_403
timestamp 1644511149
transform 1 0 38180 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_411
timestamp 1644511149
transform 1 0 38916 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_437
timestamp 1644511149
transform 1 0 41308 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_449
timestamp 1644511149
transform 1 0 42412 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_455
timestamp 1644511149
transform 1 0 42964 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_70_466
timestamp 1644511149
transform 1 0 43976 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_474
timestamp 1644511149
transform 1 0 44712 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_481
timestamp 1644511149
transform 1 0 45356 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_486
timestamp 1644511149
transform 1 0 45816 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_494
timestamp 1644511149
transform 1 0 46552 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_511
timestamp 1644511149
transform 1 0 48116 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_517
timestamp 1644511149
transform 1 0 48668 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_521
timestamp 1644511149
transform 1 0 49036 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_529
timestamp 1644511149
transform 1 0 49772 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_533
timestamp 1644511149
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_545
timestamp 1644511149
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_557
timestamp 1644511149
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_569
timestamp 1644511149
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1644511149
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1644511149
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_589
timestamp 1644511149
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_601
timestamp 1644511149
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_613
timestamp 1644511149
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_625
timestamp 1644511149
transform 1 0 58604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_637
timestamp 1644511149
transform 1 0 59708 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_643
timestamp 1644511149
transform 1 0 60260 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_645
timestamp 1644511149
transform 1 0 60444 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_657
timestamp 1644511149
transform 1 0 61548 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_669
timestamp 1644511149
transform 1 0 62652 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_681
timestamp 1644511149
transform 1 0 63756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_693
timestamp 1644511149
transform 1 0 64860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1644511149
transform 1 0 65412 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_701
timestamp 1644511149
transform 1 0 65596 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_707
timestamp 1644511149
transform 1 0 66148 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_729
timestamp 1644511149
transform 1 0 68172 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1644511149
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_180
timestamp 1644511149
transform 1 0 17664 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_192
timestamp 1644511149
transform 1 0 18768 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_198
timestamp 1644511149
transform 1 0 19320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_202
timestamp 1644511149
transform 1 0 19688 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_214
timestamp 1644511149
transform 1 0 20792 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1644511149
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_233
timestamp 1644511149
transform 1 0 22540 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_71_247
timestamp 1644511149
transform 1 0 23828 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_255
timestamp 1644511149
transform 1 0 24564 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_260
timestamp 1644511149
transform 1 0 25024 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_267
timestamp 1644511149
transform 1 0 25668 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_285
timestamp 1644511149
transform 1 0 27324 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_290
timestamp 1644511149
transform 1 0 27784 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_301
timestamp 1644511149
transform 1 0 28796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_308
timestamp 1644511149
transform 1 0 29440 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_324
timestamp 1644511149
transform 1 0 30912 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_362
timestamp 1644511149
transform 1 0 34408 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_366
timestamp 1644511149
transform 1 0 34776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_383
timestamp 1644511149
transform 1 0 36340 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_398
timestamp 1644511149
transform 1 0 37720 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_406
timestamp 1644511149
transform 1 0 38456 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_410
timestamp 1644511149
transform 1 0 38824 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_427
timestamp 1644511149
transform 1 0 40388 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_433
timestamp 1644511149
transform 1 0 40940 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_444
timestamp 1644511149
transform 1 0 41952 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_456
timestamp 1644511149
transform 1 0 43056 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_464
timestamp 1644511149
transform 1 0 43792 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_471
timestamp 1644511149
transform 1 0 44436 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_483
timestamp 1644511149
transform 1 0 45540 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_493
timestamp 1644511149
transform 1 0 46460 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_501
timestamp 1644511149
transform 1 0 47196 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_538
timestamp 1644511149
transform 1 0 50600 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_550
timestamp 1644511149
transform 1 0 51704 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_558
timestamp 1644511149
transform 1 0 52440 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_561
timestamp 1644511149
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_573
timestamp 1644511149
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_585
timestamp 1644511149
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_597
timestamp 1644511149
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1644511149
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1644511149
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_617
timestamp 1644511149
transform 1 0 57868 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_629
timestamp 1644511149
transform 1 0 58972 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_641
timestamp 1644511149
transform 1 0 60076 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_653
timestamp 1644511149
transform 1 0 61180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_665
timestamp 1644511149
transform 1 0 62284 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_671
timestamp 1644511149
transform 1 0 62836 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_673
timestamp 1644511149
transform 1 0 63020 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_685
timestamp 1644511149
transform 1 0 64124 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_697
timestamp 1644511149
transform 1 0 65228 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_709
timestamp 1644511149
transform 1 0 66332 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_713
timestamp 1644511149
transform 1 0 66700 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_717
timestamp 1644511149
transform 1 0 67068 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_724
timestamp 1644511149
transform 1 0 67712 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_729
timestamp 1644511149
transform 1 0 68172 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1644511149
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1644511149
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_160
timestamp 1644511149
transform 1 0 15824 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_174
timestamp 1644511149
transform 1 0 17112 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_183
timestamp 1644511149
transform 1 0 17940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_213
timestamp 1644511149
transform 1 0 20700 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_241
timestamp 1644511149
transform 1 0 23276 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_246
timestamp 1644511149
transform 1 0 23736 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_256
timestamp 1644511149
transform 1 0 24656 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_270
timestamp 1644511149
transform 1 0 25944 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_278
timestamp 1644511149
transform 1 0 26680 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_282
timestamp 1644511149
transform 1 0 27048 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_304
timestamp 1644511149
transform 1 0 29072 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_329
timestamp 1644511149
transform 1 0 31372 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_335
timestamp 1644511149
transform 1 0 31924 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_340
timestamp 1644511149
transform 1 0 32384 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_348
timestamp 1644511149
transform 1 0 33120 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_352
timestamp 1644511149
transform 1 0 33488 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_72_374
timestamp 1644511149
transform 1 0 35512 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_382
timestamp 1644511149
transform 1 0 36248 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_388
timestamp 1644511149
transform 1 0 36800 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_397
timestamp 1644511149
transform 1 0 37628 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_439
timestamp 1644511149
transform 1 0 41492 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_443
timestamp 1644511149
transform 1 0 41860 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_451
timestamp 1644511149
transform 1 0 42596 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_460
timestamp 1644511149
transform 1 0 43424 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_472
timestamp 1644511149
transform 1 0 44528 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_487
timestamp 1644511149
transform 1 0 45908 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_507
timestamp 1644511149
transform 1 0 47748 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_515
timestamp 1644511149
transform 1 0 48484 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_520
timestamp 1644511149
transform 1 0 48944 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_527
timestamp 1644511149
transform 1 0 49588 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1644511149
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_533
timestamp 1644511149
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_545
timestamp 1644511149
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_557
timestamp 1644511149
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_569
timestamp 1644511149
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1644511149
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1644511149
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_589
timestamp 1644511149
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_601
timestamp 1644511149
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_613
timestamp 1644511149
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_625
timestamp 1644511149
transform 1 0 58604 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_637
timestamp 1644511149
transform 1 0 59708 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_643
timestamp 1644511149
transform 1 0 60260 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_645
timestamp 1644511149
transform 1 0 60444 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_657
timestamp 1644511149
transform 1 0 61548 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_669
timestamp 1644511149
transform 1 0 62652 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_681
timestamp 1644511149
transform 1 0 63756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_693
timestamp 1644511149
transform 1 0 64860 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1644511149
transform 1 0 65412 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_701
timestamp 1644511149
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_713
timestamp 1644511149
transform 1 0 66700 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_721
timestamp 1644511149
transform 1 0 67436 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_725
timestamp 1644511149
transform 1 0 67804 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1644511149
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1644511149
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1644511149
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_145
timestamp 1644511149
transform 1 0 14444 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_164
timestamp 1644511149
transform 1 0 16192 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_188
timestamp 1644511149
transform 1 0 18400 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_196
timestamp 1644511149
transform 1 0 19136 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_235
timestamp 1644511149
transform 1 0 22724 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_243
timestamp 1644511149
transform 1 0 23460 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_251
timestamp 1644511149
transform 1 0 24196 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_257
timestamp 1644511149
transform 1 0 24748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_263
timestamp 1644511149
transform 1 0 25300 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_267
timestamp 1644511149
transform 1 0 25668 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_275
timestamp 1644511149
transform 1 0 26404 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_298
timestamp 1644511149
transform 1 0 28520 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_325
timestamp 1644511149
transform 1 0 31004 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_332
timestamp 1644511149
transform 1 0 31648 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_353
timestamp 1644511149
transform 1 0 33580 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_369
timestamp 1644511149
transform 1 0 35052 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_376
timestamp 1644511149
transform 1 0 35696 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_382
timestamp 1644511149
transform 1 0 36248 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_388
timestamp 1644511149
transform 1 0 36800 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_398
timestamp 1644511149
transform 1 0 37720 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_404
timestamp 1644511149
transform 1 0 38272 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_412
timestamp 1644511149
transform 1 0 39008 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_421
timestamp 1644511149
transform 1 0 39836 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_433
timestamp 1644511149
transform 1 0 40940 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_460
timestamp 1644511149
transform 1 0 43424 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_480
timestamp 1644511149
transform 1 0 45264 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_492
timestamp 1644511149
transform 1 0 46368 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_513
timestamp 1644511149
transform 1 0 48300 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_537
timestamp 1644511149
transform 1 0 50508 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_549
timestamp 1644511149
transform 1 0 51612 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_557
timestamp 1644511149
transform 1 0 52348 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_561
timestamp 1644511149
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_573
timestamp 1644511149
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_585
timestamp 1644511149
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_597
timestamp 1644511149
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1644511149
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1644511149
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_617
timestamp 1644511149
transform 1 0 57868 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_629
timestamp 1644511149
transform 1 0 58972 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_641
timestamp 1644511149
transform 1 0 60076 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_653
timestamp 1644511149
transform 1 0 61180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_665
timestamp 1644511149
transform 1 0 62284 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_671
timestamp 1644511149
transform 1 0 62836 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_673
timestamp 1644511149
transform 1 0 63020 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_685
timestamp 1644511149
transform 1 0 64124 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_697
timestamp 1644511149
transform 1 0 65228 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_724
timestamp 1644511149
transform 1 0 67712 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_729
timestamp 1644511149
transform 1 0 68172 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_11
timestamp 1644511149
transform 1 0 2116 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_23
timestamp 1644511149
transform 1 0 3220 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_129
timestamp 1644511149
transform 1 0 12972 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_134
timestamp 1644511149
transform 1 0 13432 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_147
timestamp 1644511149
transform 1 0 14628 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_152
timestamp 1644511149
transform 1 0 15088 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_159
timestamp 1644511149
transform 1 0 15732 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_175
timestamp 1644511149
transform 1 0 17204 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_184
timestamp 1644511149
transform 1 0 18032 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_217
timestamp 1644511149
transform 1 0 21068 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_224
timestamp 1644511149
transform 1 0 21712 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_236
timestamp 1644511149
transform 1 0 22816 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_242
timestamp 1644511149
transform 1 0 23368 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_247
timestamp 1644511149
transform 1 0 23828 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_269
timestamp 1644511149
transform 1 0 25852 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_281
timestamp 1644511149
transform 1 0 26956 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_293
timestamp 1644511149
transform 1 0 28060 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_305
timestamp 1644511149
transform 1 0 29164 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_319
timestamp 1644511149
transform 1 0 30452 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_327
timestamp 1644511149
transform 1 0 31188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_336
timestamp 1644511149
transform 1 0 32016 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_353
timestamp 1644511149
transform 1 0 33580 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_360
timestamp 1644511149
transform 1 0 34224 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_381
timestamp 1644511149
transform 1 0 36156 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_387
timestamp 1644511149
transform 1 0 36708 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_398
timestamp 1644511149
transform 1 0 37720 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_407
timestamp 1644511149
transform 1 0 38548 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_415
timestamp 1644511149
transform 1 0 39284 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_426
timestamp 1644511149
transform 1 0 40296 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_434
timestamp 1644511149
transform 1 0 41032 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_451
timestamp 1644511149
transform 1 0 42596 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_458
timestamp 1644511149
transform 1 0 43240 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_472
timestamp 1644511149
transform 1 0 44528 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_480
timestamp 1644511149
transform 1 0 45264 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_492
timestamp 1644511149
transform 1 0 46368 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_504
timestamp 1644511149
transform 1 0 47472 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_508
timestamp 1644511149
transform 1 0 47840 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_524
timestamp 1644511149
transform 1 0 49312 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_533
timestamp 1644511149
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_545
timestamp 1644511149
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_557
timestamp 1644511149
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_569
timestamp 1644511149
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1644511149
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1644511149
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_589
timestamp 1644511149
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_601
timestamp 1644511149
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_613
timestamp 1644511149
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_625
timestamp 1644511149
transform 1 0 58604 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_637
timestamp 1644511149
transform 1 0 59708 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_643
timestamp 1644511149
transform 1 0 60260 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_645
timestamp 1644511149
transform 1 0 60444 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_657
timestamp 1644511149
transform 1 0 61548 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_669
timestamp 1644511149
transform 1 0 62652 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_681
timestamp 1644511149
transform 1 0 63756 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1644511149
transform 1 0 64860 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1644511149
transform 1 0 65412 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_701
timestamp 1644511149
transform 1 0 65596 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_713
timestamp 1644511149
transform 1 0 66700 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_720
timestamp 1644511149
transform 1 0 67344 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_727
timestamp 1644511149
transform 1 0 67988 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_142
timestamp 1644511149
transform 1 0 14168 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_150
timestamp 1644511149
transform 1 0 14904 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_159
timestamp 1644511149
transform 1 0 15732 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_174
timestamp 1644511149
transform 1 0 17112 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_186
timestamp 1644511149
transform 1 0 18216 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_194
timestamp 1644511149
transform 1 0 18952 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_218
timestamp 1644511149
transform 1 0 21160 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_243
timestamp 1644511149
transform 1 0 23460 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_247
timestamp 1644511149
transform 1 0 23828 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_252
timestamp 1644511149
transform 1 0 24288 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_260
timestamp 1644511149
transform 1 0 25024 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_268
timestamp 1644511149
transform 1 0 25760 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_297
timestamp 1644511149
transform 1 0 28428 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_75_326
timestamp 1644511149
transform 1 0 31096 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_334
timestamp 1644511149
transform 1 0 31832 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_345
timestamp 1644511149
transform 1 0 32844 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_351
timestamp 1644511149
transform 1 0 33396 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_360
timestamp 1644511149
transform 1 0 34224 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_368
timestamp 1644511149
transform 1 0 34960 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_380
timestamp 1644511149
transform 1 0 36064 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_399
timestamp 1644511149
transform 1 0 37812 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_406
timestamp 1644511149
transform 1 0 38456 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_426
timestamp 1644511149
transform 1 0 40296 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_436
timestamp 1644511149
transform 1 0 41216 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_444
timestamp 1644511149
transform 1 0 41952 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_468
timestamp 1644511149
transform 1 0 44160 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_480
timestamp 1644511149
transform 1 0 45264 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_488
timestamp 1644511149
transform 1 0 46000 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_495
timestamp 1644511149
transform 1 0 46644 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1644511149
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_510
timestamp 1644511149
transform 1 0 48024 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_518
timestamp 1644511149
transform 1 0 48760 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_530
timestamp 1644511149
transform 1 0 49864 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_542
timestamp 1644511149
transform 1 0 50968 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_554
timestamp 1644511149
transform 1 0 52072 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_561
timestamp 1644511149
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_573
timestamp 1644511149
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_585
timestamp 1644511149
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_597
timestamp 1644511149
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1644511149
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1644511149
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_617
timestamp 1644511149
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_629
timestamp 1644511149
transform 1 0 58972 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_641
timestamp 1644511149
transform 1 0 60076 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_653
timestamp 1644511149
transform 1 0 61180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_665
timestamp 1644511149
transform 1 0 62284 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_671
timestamp 1644511149
transform 1 0 62836 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_673
timestamp 1644511149
transform 1 0 63020 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_685
timestamp 1644511149
transform 1 0 64124 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_697
timestamp 1644511149
transform 1 0 65228 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_709
timestamp 1644511149
transform 1 0 66332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_724
timestamp 1644511149
transform 1 0 67712 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_729
timestamp 1644511149
transform 1 0 68172 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_11
timestamp 1644511149
transform 1 0 2116 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_23
timestamp 1644511149
transform 1 0 3220 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_129
timestamp 1644511149
transform 1 0 12972 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_136
timestamp 1644511149
transform 1 0 13616 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_76_163
timestamp 1644511149
transform 1 0 16100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_169
timestamp 1644511149
transform 1 0 16652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_186
timestamp 1644511149
transform 1 0 18216 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_194
timestamp 1644511149
transform 1 0 18952 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_205
timestamp 1644511149
transform 1 0 19964 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_211
timestamp 1644511149
transform 1 0 20516 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_231
timestamp 1644511149
transform 1 0 22356 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_269
timestamp 1644511149
transform 1 0 25852 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_304
timestamp 1644511149
transform 1 0 29072 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_314
timestamp 1644511149
transform 1 0 29992 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_322
timestamp 1644511149
transform 1 0 30728 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_340
timestamp 1644511149
transform 1 0 32384 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_360
timestamp 1644511149
transform 1 0 34224 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_386
timestamp 1644511149
transform 1 0 36616 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_398
timestamp 1644511149
transform 1 0 37720 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_404
timestamp 1644511149
transform 1 0 38272 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_427
timestamp 1644511149
transform 1 0 40388 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_435
timestamp 1644511149
transform 1 0 41124 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_447
timestamp 1644511149
transform 1 0 42228 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_452
timestamp 1644511149
transform 1 0 42688 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_464
timestamp 1644511149
transform 1 0 43792 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_471
timestamp 1644511149
transform 1 0 44436 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_500
timestamp 1644511149
transform 1 0 47104 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_508
timestamp 1644511149
transform 1 0 47840 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_526
timestamp 1644511149
transform 1 0 49496 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_533
timestamp 1644511149
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_545
timestamp 1644511149
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_557
timestamp 1644511149
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_569
timestamp 1644511149
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1644511149
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1644511149
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_589
timestamp 1644511149
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_601
timestamp 1644511149
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_613
timestamp 1644511149
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_625
timestamp 1644511149
transform 1 0 58604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_637
timestamp 1644511149
transform 1 0 59708 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_643
timestamp 1644511149
transform 1 0 60260 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_645
timestamp 1644511149
transform 1 0 60444 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_657
timestamp 1644511149
transform 1 0 61548 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_669
timestamp 1644511149
transform 1 0 62652 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_681
timestamp 1644511149
transform 1 0 63756 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_693
timestamp 1644511149
transform 1 0 64860 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_699
timestamp 1644511149
transform 1 0 65412 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_701
timestamp 1644511149
transform 1 0 65596 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_707
timestamp 1644511149
transform 1 0 66148 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_729
timestamp 1644511149
transform 1 0 68172 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_129
timestamp 1644511149
transform 1 0 12972 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_141
timestamp 1644511149
transform 1 0 14076 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_156
timestamp 1644511149
transform 1 0 15456 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_172
timestamp 1644511149
transform 1 0 16928 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_180
timestamp 1644511149
transform 1 0 17664 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_204
timestamp 1644511149
transform 1 0 19872 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_216
timestamp 1644511149
transform 1 0 20976 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_244
timestamp 1644511149
transform 1 0 23552 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_256
timestamp 1644511149
transform 1 0 24656 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_263
timestamp 1644511149
transform 1 0 25300 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_275
timestamp 1644511149
transform 1 0 26404 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_284
timestamp 1644511149
transform 1 0 27232 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_296
timestamp 1644511149
transform 1 0 28336 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_308
timestamp 1644511149
transform 1 0 29440 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_318
timestamp 1644511149
transform 1 0 30360 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_327
timestamp 1644511149
transform 1 0 31188 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_340
timestamp 1644511149
transform 1 0 32384 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_352
timestamp 1644511149
transform 1 0 33488 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_77_358
timestamp 1644511149
transform 1 0 34040 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_368
timestamp 1644511149
transform 1 0 34960 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_388
timestamp 1644511149
transform 1 0 36800 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_437
timestamp 1644511149
transform 1 0 41308 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_444
timestamp 1644511149
transform 1 0 41952 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_453
timestamp 1644511149
transform 1 0 42780 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_481
timestamp 1644511149
transform 1 0 45356 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_487
timestamp 1644511149
transform 1 0 45908 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_494
timestamp 1644511149
transform 1 0 46552 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_502
timestamp 1644511149
transform 1 0 47288 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_510
timestamp 1644511149
transform 1 0 48024 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_518
timestamp 1644511149
transform 1 0 48760 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_522
timestamp 1644511149
transform 1 0 49128 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_527
timestamp 1644511149
transform 1 0 49588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_539
timestamp 1644511149
transform 1 0 50692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_551
timestamp 1644511149
transform 1 0 51796 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1644511149
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_561
timestamp 1644511149
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_573
timestamp 1644511149
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_585
timestamp 1644511149
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_597
timestamp 1644511149
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1644511149
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1644511149
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_617
timestamp 1644511149
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_629
timestamp 1644511149
transform 1 0 58972 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_641
timestamp 1644511149
transform 1 0 60076 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_653
timestamp 1644511149
transform 1 0 61180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1644511149
transform 1 0 62284 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1644511149
transform 1 0 62836 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_673
timestamp 1644511149
transform 1 0 63020 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_685
timestamp 1644511149
transform 1 0 64124 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_697
timestamp 1644511149
transform 1 0 65228 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_709
timestamp 1644511149
transform 1 0 66332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_724
timestamp 1644511149
transform 1 0 67712 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_729
timestamp 1644511149
transform 1 0 68172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_127
timestamp 1644511149
transform 1 0 12788 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_136
timestamp 1644511149
transform 1 0 13616 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_149
timestamp 1644511149
transform 1 0 14812 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_157
timestamp 1644511149
transform 1 0 15548 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_169
timestamp 1644511149
transform 1 0 16652 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_181
timestamp 1644511149
transform 1 0 17756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_193
timestamp 1644511149
transform 1 0 18860 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_201
timestamp 1644511149
transform 1 0 19596 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_208
timestamp 1644511149
transform 1 0 20240 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_220
timestamp 1644511149
transform 1 0 21344 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_227
timestamp 1644511149
transform 1 0 21988 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_235
timestamp 1644511149
transform 1 0 22724 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_78_241
timestamp 1644511149
transform 1 0 23276 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_249
timestamp 1644511149
transform 1 0 24012 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_271
timestamp 1644511149
transform 1 0 26036 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_283
timestamp 1644511149
transform 1 0 27140 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_78_290
timestamp 1644511149
transform 1 0 27784 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_298
timestamp 1644511149
transform 1 0 28520 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_304
timestamp 1644511149
transform 1 0 29072 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_315
timestamp 1644511149
transform 1 0 30084 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_320
timestamp 1644511149
transform 1 0 30544 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_328
timestamp 1644511149
transform 1 0 31280 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_340
timestamp 1644511149
transform 1 0 32384 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_344
timestamp 1644511149
transform 1 0 32752 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_356
timestamp 1644511149
transform 1 0 33856 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_383
timestamp 1644511149
transform 1 0 36340 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_398
timestamp 1644511149
transform 1 0 37720 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_407
timestamp 1644511149
transform 1 0 38548 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_426
timestamp 1644511149
transform 1 0 40296 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_438
timestamp 1644511149
transform 1 0 41400 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_78_457
timestamp 1644511149
transform 1 0 43148 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_463
timestamp 1644511149
transform 1 0 43700 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_467
timestamp 1644511149
transform 1 0 44068 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1644511149
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_485
timestamp 1644511149
transform 1 0 45724 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_501
timestamp 1644511149
transform 1 0 47196 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_521
timestamp 1644511149
transform 1 0 49036 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_529
timestamp 1644511149
transform 1 0 49772 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_537
timestamp 1644511149
transform 1 0 50508 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_549
timestamp 1644511149
transform 1 0 51612 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_561
timestamp 1644511149
transform 1 0 52716 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_573
timestamp 1644511149
transform 1 0 53820 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_585
timestamp 1644511149
transform 1 0 54924 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_589
timestamp 1644511149
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_601
timestamp 1644511149
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_613
timestamp 1644511149
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_625
timestamp 1644511149
transform 1 0 58604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1644511149
transform 1 0 59708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1644511149
transform 1 0 60260 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_645
timestamp 1644511149
transform 1 0 60444 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_657
timestamp 1644511149
transform 1 0 61548 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_669
timestamp 1644511149
transform 1 0 62652 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_681
timestamp 1644511149
transform 1 0 63756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_693
timestamp 1644511149
transform 1 0 64860 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_699
timestamp 1644511149
transform 1 0 65412 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_701
timestamp 1644511149
transform 1 0 65596 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_707
timestamp 1644511149
transform 1 0 66148 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_729
timestamp 1644511149
transform 1 0 68172 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_11
timestamp 1644511149
transform 1 0 2116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_23
timestamp 1644511149
transform 1 0 3220 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_35
timestamp 1644511149
transform 1 0 4324 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_47
timestamp 1644511149
transform 1 0 5428 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_121
timestamp 1644511149
transform 1 0 12236 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_79_140
timestamp 1644511149
transform 1 0 13984 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_79_162
timestamp 1644511149
transform 1 0 16008 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_173
timestamp 1644511149
transform 1 0 17020 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_177
timestamp 1644511149
transform 1 0 17388 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_199
timestamp 1644511149
transform 1 0 19412 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_219
timestamp 1644511149
transform 1 0 21252 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_231
timestamp 1644511149
transform 1 0 22356 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_239
timestamp 1644511149
transform 1 0 23092 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_257
timestamp 1644511149
transform 1 0 24748 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_265
timestamp 1644511149
transform 1 0 25484 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_271
timestamp 1644511149
transform 1 0 26036 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_284
timestamp 1644511149
transform 1 0 27232 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_304
timestamp 1644511149
transform 1 0 29072 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_313
timestamp 1644511149
transform 1 0 29900 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_323
timestamp 1644511149
transform 1 0 30820 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_79_348
timestamp 1644511149
transform 1 0 33120 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_356
timestamp 1644511149
transform 1 0 33856 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_369
timestamp 1644511149
transform 1 0 35052 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_376
timestamp 1644511149
transform 1 0 35696 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_388
timestamp 1644511149
transform 1 0 36800 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_409
timestamp 1644511149
transform 1 0 38732 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_437
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_445
timestamp 1644511149
transform 1 0 42044 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_453
timestamp 1644511149
transform 1 0 42780 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_465
timestamp 1644511149
transform 1 0 43884 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_473
timestamp 1644511149
transform 1 0 44620 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_482
timestamp 1644511149
transform 1 0 45448 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_494
timestamp 1644511149
transform 1 0 46552 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_502
timestamp 1644511149
transform 1 0 47288 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_509
timestamp 1644511149
transform 1 0 47932 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_516
timestamp 1644511149
transform 1 0 48576 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_528
timestamp 1644511149
transform 1 0 49680 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_532
timestamp 1644511149
transform 1 0 50048 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_549
timestamp 1644511149
transform 1 0 51612 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_557
timestamp 1644511149
transform 1 0 52348 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_561
timestamp 1644511149
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_573
timestamp 1644511149
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_585
timestamp 1644511149
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_597
timestamp 1644511149
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1644511149
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1644511149
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_617
timestamp 1644511149
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_629
timestamp 1644511149
transform 1 0 58972 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_641
timestamp 1644511149
transform 1 0 60076 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_653
timestamp 1644511149
transform 1 0 61180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_665
timestamp 1644511149
transform 1 0 62284 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_671
timestamp 1644511149
transform 1 0 62836 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_673
timestamp 1644511149
transform 1 0 63020 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_685
timestamp 1644511149
transform 1 0 64124 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_697
timestamp 1644511149
transform 1 0 65228 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_709
timestamp 1644511149
transform 1 0 66332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_724
timestamp 1644511149
transform 1 0 67712 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_729
timestamp 1644511149
transform 1 0 68172 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_80_132
timestamp 1644511149
transform 1 0 13248 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_149
timestamp 1644511149
transform 1 0 14812 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_156
timestamp 1644511149
transform 1 0 15456 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_164
timestamp 1644511149
transform 1 0 16192 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_183
timestamp 1644511149
transform 1 0 17940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_190
timestamp 1644511149
transform 1 0 18584 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_201
timestamp 1644511149
transform 1 0 19596 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_207
timestamp 1644511149
transform 1 0 20148 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_216
timestamp 1644511149
transform 1 0 20976 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_222
timestamp 1644511149
transform 1 0 21528 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_239
timestamp 1644511149
transform 1 0 23092 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_248
timestamp 1644511149
transform 1 0 23920 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_258
timestamp 1644511149
transform 1 0 24840 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_266
timestamp 1644511149
transform 1 0 25576 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_284
timestamp 1644511149
transform 1 0 27232 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_299
timestamp 1644511149
transform 1 0 28612 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_329
timestamp 1644511149
transform 1 0 31372 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_335
timestamp 1644511149
transform 1 0 31924 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_352
timestamp 1644511149
transform 1 0 33488 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_359
timestamp 1644511149
transform 1 0 34132 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_372
timestamp 1644511149
transform 1 0 35328 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_382
timestamp 1644511149
transform 1 0 36248 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_390
timestamp 1644511149
transform 1 0 36984 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_402
timestamp 1644511149
transform 1 0 38088 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_414
timestamp 1644511149
transform 1 0 39192 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_439
timestamp 1644511149
transform 1 0 41492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_461
timestamp 1644511149
transform 1 0 43516 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_473
timestamp 1644511149
transform 1 0 44620 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_481
timestamp 1644511149
transform 1 0 45356 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_488
timestamp 1644511149
transform 1 0 46000 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_500
timestamp 1644511149
transform 1 0 47104 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_508
timestamp 1644511149
transform 1 0 47840 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_514
timestamp 1644511149
transform 1 0 48392 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_526
timestamp 1644511149
transform 1 0 49496 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_533
timestamp 1644511149
transform 1 0 50140 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_537
timestamp 1644511149
transform 1 0 50508 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_543
timestamp 1644511149
transform 1 0 51060 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_550
timestamp 1644511149
transform 1 0 51704 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_562
timestamp 1644511149
transform 1 0 52808 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_574
timestamp 1644511149
transform 1 0 53912 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_586
timestamp 1644511149
transform 1 0 55016 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_589
timestamp 1644511149
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_601
timestamp 1644511149
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_613
timestamp 1644511149
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_625
timestamp 1644511149
transform 1 0 58604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_637
timestamp 1644511149
transform 1 0 59708 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_643
timestamp 1644511149
transform 1 0 60260 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_645
timestamp 1644511149
transform 1 0 60444 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_657
timestamp 1644511149
transform 1 0 61548 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_669
timestamp 1644511149
transform 1 0 62652 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_681
timestamp 1644511149
transform 1 0 63756 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_693
timestamp 1644511149
transform 1 0 64860 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_699
timestamp 1644511149
transform 1 0 65412 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_701
timestamp 1644511149
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_713
timestamp 1644511149
transform 1 0 66700 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_80_722
timestamp 1644511149
transform 1 0 67528 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_730
timestamp 1644511149
transform 1 0 68264 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_11
timestamp 1644511149
transform 1 0 2116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_23
timestamp 1644511149
transform 1 0 3220 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_35
timestamp 1644511149
transform 1 0 4324 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_47
timestamp 1644511149
transform 1 0 5428 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_175
timestamp 1644511149
transform 1 0 17204 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_199
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_203
timestamp 1644511149
transform 1 0 19780 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_229
timestamp 1644511149
transform 1 0 22172 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_236
timestamp 1644511149
transform 1 0 22816 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_248
timestamp 1644511149
transform 1 0 23920 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_270
timestamp 1644511149
transform 1 0 25944 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1644511149
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_301
timestamp 1644511149
transform 1 0 28796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_310
timestamp 1644511149
transform 1 0 29624 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_318
timestamp 1644511149
transform 1 0 30360 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_325
timestamp 1644511149
transform 1 0 31004 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_333
timestamp 1644511149
transform 1 0 31740 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_343
timestamp 1644511149
transform 1 0 32660 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_354
timestamp 1644511149
transform 1 0 33672 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_378
timestamp 1644511149
transform 1 0 35880 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_386
timestamp 1644511149
transform 1 0 36616 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_403
timestamp 1644511149
transform 1 0 38180 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_411
timestamp 1644511149
transform 1 0 38916 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_415
timestamp 1644511149
transform 1 0 39284 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_420
timestamp 1644511149
transform 1 0 39744 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_432
timestamp 1644511149
transform 1 0 40848 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_440
timestamp 1644511149
transform 1 0 41584 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1644511149
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_453
timestamp 1644511149
transform 1 0 42780 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_464
timestamp 1644511149
transform 1 0 43792 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_487
timestamp 1644511149
transform 1 0 45908 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_495
timestamp 1644511149
transform 1 0 46644 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_521
timestamp 1644511149
transform 1 0 49036 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_541
timestamp 1644511149
transform 1 0 50876 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_547
timestamp 1644511149
transform 1 0 51428 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1644511149
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1644511149
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_561
timestamp 1644511149
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_573
timestamp 1644511149
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_585
timestamp 1644511149
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_597
timestamp 1644511149
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1644511149
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1644511149
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_617
timestamp 1644511149
transform 1 0 57868 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_629
timestamp 1644511149
transform 1 0 58972 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_641
timestamp 1644511149
transform 1 0 60076 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_653
timestamp 1644511149
transform 1 0 61180 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_665
timestamp 1644511149
transform 1 0 62284 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_671
timestamp 1644511149
transform 1 0 62836 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_673
timestamp 1644511149
transform 1 0 63020 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_685
timestamp 1644511149
transform 1 0 64124 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_697
timestamp 1644511149
transform 1 0 65228 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_724
timestamp 1644511149
transform 1 0 67712 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_729
timestamp 1644511149
transform 1 0 68172 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_11
timestamp 1644511149
transform 1 0 2116 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_16
timestamp 1644511149
transform 1 0 2576 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1644511149
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_65
timestamp 1644511149
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1644511149
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_134
timestamp 1644511149
transform 1 0 13432 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_149
timestamp 1644511149
transform 1 0 14812 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_155
timestamp 1644511149
transform 1 0 15364 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_163
timestamp 1644511149
transform 1 0 16100 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_181
timestamp 1644511149
transform 1 0 17756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_193
timestamp 1644511149
transform 1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_205
timestamp 1644511149
transform 1 0 19964 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_210
timestamp 1644511149
transform 1 0 20424 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_217
timestamp 1644511149
transform 1 0 21068 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_235
timestamp 1644511149
transform 1 0 22724 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_242
timestamp 1644511149
transform 1 0 23368 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1644511149
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_273
timestamp 1644511149
transform 1 0 26220 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_291
timestamp 1644511149
transform 1 0 27876 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_299
timestamp 1644511149
transform 1 0 28612 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_304
timestamp 1644511149
transform 1 0 29072 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_314
timestamp 1644511149
transform 1 0 29992 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_329
timestamp 1644511149
transform 1 0 31372 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_336
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_344
timestamp 1644511149
transform 1 0 32752 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_352
timestamp 1644511149
transform 1 0 33488 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_360
timestamp 1644511149
transform 1 0 34224 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_369
timestamp 1644511149
transform 1 0 35052 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_390
timestamp 1644511149
transform 1 0 36984 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1644511149
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1644511149
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_426
timestamp 1644511149
transform 1 0 40296 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_437
timestamp 1644511149
transform 1 0 41308 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_461
timestamp 1644511149
transform 1 0 43516 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1644511149
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1644511149
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_487
timestamp 1644511149
transform 1 0 45908 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_496
timestamp 1644511149
transform 1 0 46736 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_508
timestamp 1644511149
transform 1 0 47840 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_520
timestamp 1644511149
transform 1 0 48944 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_533
timestamp 1644511149
transform 1 0 50140 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_545
timestamp 1644511149
transform 1 0 51244 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_565
timestamp 1644511149
transform 1 0 53084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_577
timestamp 1644511149
transform 1 0 54188 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_585
timestamp 1644511149
transform 1 0 54924 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_589
timestamp 1644511149
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_601
timestamp 1644511149
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_613
timestamp 1644511149
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_625
timestamp 1644511149
transform 1 0 58604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_637
timestamp 1644511149
transform 1 0 59708 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_643
timestamp 1644511149
transform 1 0 60260 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_645
timestamp 1644511149
transform 1 0 60444 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_657
timestamp 1644511149
transform 1 0 61548 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_669
timestamp 1644511149
transform 1 0 62652 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_681
timestamp 1644511149
transform 1 0 63756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_693
timestamp 1644511149
transform 1 0 64860 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_699
timestamp 1644511149
transform 1 0 65412 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_701
timestamp 1644511149
transform 1 0 65596 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_713
timestamp 1644511149
transform 1 0 66700 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_721
timestamp 1644511149
transform 1 0 67436 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_82_727
timestamp 1644511149
transform 1 0 67988 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_83_3
timestamp 1644511149
transform 1 0 1380 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_27
timestamp 1644511149
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_39
timestamp 1644511149
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1644511149
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1644511149
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1644511149
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1644511149
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_81
timestamp 1644511149
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_93
timestamp 1644511149
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1644511149
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1644511149
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_113
timestamp 1644511149
transform 1 0 11500 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_119
timestamp 1644511149
transform 1 0 12052 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_136
timestamp 1644511149
transform 1 0 13616 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_83_158
timestamp 1644511149
transform 1 0 15640 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_166
timestamp 1644511149
transform 1 0 16376 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_169
timestamp 1644511149
transform 1 0 16652 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_178
timestamp 1644511149
transform 1 0 17480 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_203
timestamp 1644511149
transform 1 0 19780 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_215
timestamp 1644511149
transform 1 0 20884 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1644511149
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_225
timestamp 1644511149
transform 1 0 21804 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_229
timestamp 1644511149
transform 1 0 22172 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_246
timestamp 1644511149
transform 1 0 23736 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_254
timestamp 1644511149
transform 1 0 24472 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_266
timestamp 1644511149
transform 1 0 25576 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_276
timestamp 1644511149
transform 1 0 26496 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_281
timestamp 1644511149
transform 1 0 26956 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_288
timestamp 1644511149
transform 1 0 27600 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_310
timestamp 1644511149
transform 1 0 29624 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_332
timestamp 1644511149
transform 1 0 31648 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_337
timestamp 1644511149
transform 1 0 32108 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_341
timestamp 1644511149
transform 1 0 32476 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_359
timestamp 1644511149
transform 1 0 34132 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_363
timestamp 1644511149
transform 1 0 34500 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_370
timestamp 1644511149
transform 1 0 35144 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_381
timestamp 1644511149
transform 1 0 36156 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_389
timestamp 1644511149
transform 1 0 36892 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_83_393
timestamp 1644511149
transform 1 0 37260 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_83_403
timestamp 1644511149
transform 1 0 38180 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_426
timestamp 1644511149
transform 1 0 40296 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_434
timestamp 1644511149
transform 1 0 41032 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1644511149
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1644511149
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_449
timestamp 1644511149
transform 1 0 42412 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_457
timestamp 1644511149
transform 1 0 43148 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_466
timestamp 1644511149
transform 1 0 43976 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_474
timestamp 1644511149
transform 1 0 44712 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_482
timestamp 1644511149
transform 1 0 45448 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_494
timestamp 1644511149
transform 1 0 46552 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_502
timestamp 1644511149
transform 1 0 47288 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_505
timestamp 1644511149
transform 1 0 47564 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_518
timestamp 1644511149
transform 1 0 48760 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_530
timestamp 1644511149
transform 1 0 49864 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_83_540
timestamp 1644511149
transform 1 0 50784 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_546
timestamp 1644511149
transform 1 0 51336 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_550
timestamp 1644511149
transform 1 0 51704 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_558
timestamp 1644511149
transform 1 0 52440 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_561
timestamp 1644511149
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_573
timestamp 1644511149
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_585
timestamp 1644511149
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_597
timestamp 1644511149
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1644511149
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1644511149
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_617
timestamp 1644511149
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_629
timestamp 1644511149
transform 1 0 58972 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_641
timestamp 1644511149
transform 1 0 60076 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_653
timestamp 1644511149
transform 1 0 61180 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_665
timestamp 1644511149
transform 1 0 62284 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_671
timestamp 1644511149
transform 1 0 62836 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_673
timestamp 1644511149
transform 1 0 63020 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_685
timestamp 1644511149
transform 1 0 64124 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_697
timestamp 1644511149
transform 1 0 65228 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_709
timestamp 1644511149
transform 1 0 66332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_721
timestamp 1644511149
transform 1 0 67436 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_727
timestamp 1644511149
transform 1 0 67988 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_729
timestamp 1644511149
transform 1 0 68172 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_3
timestamp 1644511149
transform 1 0 1380 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_10
timestamp 1644511149
transform 1 0 2024 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_22
timestamp 1644511149
transform 1 0 3128 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1644511149
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1644511149
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1644511149
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1644511149
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1644511149
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1644511149
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_85
timestamp 1644511149
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_97
timestamp 1644511149
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_109
timestamp 1644511149
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_121
timestamp 1644511149
transform 1 0 12236 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_125
timestamp 1644511149
transform 1 0 12604 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_129
timestamp 1644511149
transform 1 0 12972 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_137
timestamp 1644511149
transform 1 0 13708 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_84_141
timestamp 1644511149
transform 1 0 14076 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_147
timestamp 1644511149
transform 1 0 14628 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_154
timestamp 1644511149
transform 1 0 15272 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_161
timestamp 1644511149
transform 1 0 15916 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_169
timestamp 1644511149
transform 1 0 16652 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_176
timestamp 1644511149
transform 1 0 17296 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_188
timestamp 1644511149
transform 1 0 18400 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_197
timestamp 1644511149
transform 1 0 19228 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_206
timestamp 1644511149
transform 1 0 20056 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_226
timestamp 1644511149
transform 1 0 21896 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_238
timestamp 1644511149
transform 1 0 23000 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_244
timestamp 1644511149
transform 1 0 23552 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_269
timestamp 1644511149
transform 1 0 25852 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_279
timestamp 1644511149
transform 1 0 26772 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_286
timestamp 1644511149
transform 1 0 27416 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_298
timestamp 1644511149
transform 1 0 28520 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_306
timestamp 1644511149
transform 1 0 29256 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_309
timestamp 1644511149
transform 1 0 29532 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_314
timestamp 1644511149
transform 1 0 29992 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_322
timestamp 1644511149
transform 1 0 30728 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_329
timestamp 1644511149
transform 1 0 31372 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_84_339
timestamp 1644511149
transform 1 0 32292 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_349
timestamp 1644511149
transform 1 0 33212 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1644511149
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1644511149
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_365
timestamp 1644511149
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_377
timestamp 1644511149
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_389
timestamp 1644511149
transform 1 0 36892 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_395
timestamp 1644511149
transform 1 0 37444 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_407
timestamp 1644511149
transform 1 0 38548 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1644511149
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_427
timestamp 1644511149
transform 1 0 40388 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_435
timestamp 1644511149
transform 1 0 41124 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_443
timestamp 1644511149
transform 1 0 41860 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_465
timestamp 1644511149
transform 1 0 43884 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_472
timestamp 1644511149
transform 1 0 44528 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_84_477
timestamp 1644511149
transform 1 0 44988 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_84_487
timestamp 1644511149
transform 1 0 45908 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_495
timestamp 1644511149
transform 1 0 46644 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_84_502
timestamp 1644511149
transform 1 0 47288 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_510
timestamp 1644511149
transform 1 0 48024 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_519
timestamp 1644511149
transform 1 0 48852 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_527
timestamp 1644511149
transform 1 0 49588 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1644511149
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_549
timestamp 1644511149
transform 1 0 51612 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_561
timestamp 1644511149
transform 1 0 52716 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_573
timestamp 1644511149
transform 1 0 53820 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_585
timestamp 1644511149
transform 1 0 54924 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_589
timestamp 1644511149
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_601
timestamp 1644511149
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_613
timestamp 1644511149
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_625
timestamp 1644511149
transform 1 0 58604 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_637
timestamp 1644511149
transform 1 0 59708 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_643
timestamp 1644511149
transform 1 0 60260 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_645
timestamp 1644511149
transform 1 0 60444 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_657
timestamp 1644511149
transform 1 0 61548 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_669
timestamp 1644511149
transform 1 0 62652 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_681
timestamp 1644511149
transform 1 0 63756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_693
timestamp 1644511149
transform 1 0 64860 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_699
timestamp 1644511149
transform 1 0 65412 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_701
timestamp 1644511149
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_713
timestamp 1644511149
transform 1 0 66700 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_721
timestamp 1644511149
transform 1 0 67436 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_729
timestamp 1644511149
transform 1 0 68172 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1644511149
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1644511149
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1644511149
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1644511149
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1644511149
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1644511149
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1644511149
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_69
timestamp 1644511149
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_81
timestamp 1644511149
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_93
timestamp 1644511149
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1644511149
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1644511149
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_113
timestamp 1644511149
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_125
timestamp 1644511149
transform 1 0 12604 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_132
timestamp 1644511149
transform 1 0 13248 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_144
timestamp 1644511149
transform 1 0 14352 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_156
timestamp 1644511149
transform 1 0 15456 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_169
timestamp 1644511149
transform 1 0 16652 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_177
timestamp 1644511149
transform 1 0 17388 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_189
timestamp 1644511149
transform 1 0 18492 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_204
timestamp 1644511149
transform 1 0 19872 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_212
timestamp 1644511149
transform 1 0 20608 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_220
timestamp 1644511149
transform 1 0 21344 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_225
timestamp 1644511149
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_237
timestamp 1644511149
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_249
timestamp 1644511149
transform 1 0 24012 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_260
timestamp 1644511149
transform 1 0 25024 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_267
timestamp 1644511149
transform 1 0 25668 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_276
timestamp 1644511149
transform 1 0 26496 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_286
timestamp 1644511149
transform 1 0 27416 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_298
timestamp 1644511149
transform 1 0 28520 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_302
timestamp 1644511149
transform 1 0 28888 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_309
timestamp 1644511149
transform 1 0 29532 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_319
timestamp 1644511149
transform 1 0 30452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_331
timestamp 1644511149
transform 1 0 31556 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1644511149
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_337
timestamp 1644511149
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_349
timestamp 1644511149
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_361
timestamp 1644511149
transform 1 0 34316 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_367
timestamp 1644511149
transform 1 0 34868 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_379
timestamp 1644511149
transform 1 0 35972 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_388
timestamp 1644511149
transform 1 0 36800 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_410
timestamp 1644511149
transform 1 0 38824 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_418
timestamp 1644511149
transform 1 0 39560 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_425
timestamp 1644511149
transform 1 0 40204 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_433
timestamp 1644511149
transform 1 0 40940 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_442
timestamp 1644511149
transform 1 0 41768 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_449
timestamp 1644511149
transform 1 0 42412 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_459
timestamp 1644511149
transform 1 0 43332 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_466
timestamp 1644511149
transform 1 0 43976 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_478
timestamp 1644511149
transform 1 0 45080 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_491
timestamp 1644511149
transform 1 0 46276 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_495
timestamp 1644511149
transform 1 0 46644 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_500
timestamp 1644511149
transform 1 0 47104 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_510
timestamp 1644511149
transform 1 0 48024 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_518
timestamp 1644511149
transform 1 0 48760 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_522
timestamp 1644511149
transform 1 0 49128 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_530
timestamp 1644511149
transform 1 0 49864 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_538
timestamp 1644511149
transform 1 0 50600 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_546
timestamp 1644511149
transform 1 0 51336 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_551
timestamp 1644511149
transform 1 0 51796 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1644511149
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_561
timestamp 1644511149
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_573
timestamp 1644511149
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_585
timestamp 1644511149
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_597
timestamp 1644511149
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1644511149
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1644511149
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_617
timestamp 1644511149
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_629
timestamp 1644511149
transform 1 0 58972 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_641
timestamp 1644511149
transform 1 0 60076 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_653
timestamp 1644511149
transform 1 0 61180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_665
timestamp 1644511149
transform 1 0 62284 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_671
timestamp 1644511149
transform 1 0 62836 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_673
timestamp 1644511149
transform 1 0 63020 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_685
timestamp 1644511149
transform 1 0 64124 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_697
timestamp 1644511149
transform 1 0 65228 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_709
timestamp 1644511149
transform 1 0 66332 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_721
timestamp 1644511149
transform 1 0 67436 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_727
timestamp 1644511149
transform 1 0 67988 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_729
timestamp 1644511149
transform 1 0 68172 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_3
timestamp 1644511149
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_15
timestamp 1644511149
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1644511149
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_29
timestamp 1644511149
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_41
timestamp 1644511149
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_53
timestamp 1644511149
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_65
timestamp 1644511149
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1644511149
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1644511149
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_85
timestamp 1644511149
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_97
timestamp 1644511149
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_109
timestamp 1644511149
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_121
timestamp 1644511149
transform 1 0 12236 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_129
timestamp 1644511149
transform 1 0 12972 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_135
timestamp 1644511149
transform 1 0 13524 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1644511149
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_86_141
timestamp 1644511149
transform 1 0 14076 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_147
timestamp 1644511149
transform 1 0 14628 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_161
timestamp 1644511149
transform 1 0 15916 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_181
timestamp 1644511149
transform 1 0 17756 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_190
timestamp 1644511149
transform 1 0 18584 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_200
timestamp 1644511149
transform 1 0 19504 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_214
timestamp 1644511149
transform 1 0 20792 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_222
timestamp 1644511149
transform 1 0 21528 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_239
timestamp 1644511149
transform 1 0 23092 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1644511149
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_253
timestamp 1644511149
transform 1 0 24380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_257
timestamp 1644511149
transform 1 0 24748 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_261
timestamp 1644511149
transform 1 0 25116 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_281
timestamp 1644511149
transform 1 0 26956 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_287
timestamp 1644511149
transform 1 0 27508 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_304
timestamp 1644511149
transform 1 0 29072 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_309
timestamp 1644511149
transform 1 0 29532 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_315
timestamp 1644511149
transform 1 0 30084 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_322
timestamp 1644511149
transform 1 0 30728 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_329
timestamp 1644511149
transform 1 0 31372 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_347
timestamp 1644511149
transform 1 0 33028 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_351
timestamp 1644511149
transform 1 0 33396 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_356
timestamp 1644511149
transform 1 0 33856 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_86_381
timestamp 1644511149
transform 1 0 36156 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_389
timestamp 1644511149
transform 1 0 36892 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_86_395
timestamp 1644511149
transform 1 0 37444 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_403
timestamp 1644511149
transform 1 0 38180 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_407
timestamp 1644511149
transform 1 0 38548 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_415
timestamp 1644511149
transform 1 0 39284 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1644511149
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_434
timestamp 1644511149
transform 1 0 41032 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_445
timestamp 1644511149
transform 1 0 42044 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_453
timestamp 1644511149
transform 1 0 42780 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_466
timestamp 1644511149
transform 1 0 43976 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_474
timestamp 1644511149
transform 1 0 44712 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_485
timestamp 1644511149
transform 1 0 45724 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_496
timestamp 1644511149
transform 1 0 46736 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_508
timestamp 1644511149
transform 1 0 47840 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_516
timestamp 1644511149
transform 1 0 48576 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_520
timestamp 1644511149
transform 1 0 48944 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_527
timestamp 1644511149
transform 1 0 49588 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1644511149
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_533
timestamp 1644511149
transform 1 0 50140 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_86_546
timestamp 1644511149
transform 1 0 51336 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_566
timestamp 1644511149
transform 1 0 53176 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_578
timestamp 1644511149
transform 1 0 54280 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_586
timestamp 1644511149
transform 1 0 55016 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_86_589
timestamp 1644511149
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_601
timestamp 1644511149
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_613
timestamp 1644511149
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_625
timestamp 1644511149
transform 1 0 58604 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_637
timestamp 1644511149
transform 1 0 59708 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_643
timestamp 1644511149
transform 1 0 60260 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_645
timestamp 1644511149
transform 1 0 60444 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_657
timestamp 1644511149
transform 1 0 61548 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_669
timestamp 1644511149
transform 1 0 62652 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_681
timestamp 1644511149
transform 1 0 63756 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_693
timestamp 1644511149
transform 1 0 64860 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_699
timestamp 1644511149
transform 1 0 65412 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_701
timestamp 1644511149
transform 1 0 65596 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_713
timestamp 1644511149
transform 1 0 66700 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_725
timestamp 1644511149
transform 1 0 67804 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1644511149
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1644511149
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1644511149
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_39
timestamp 1644511149
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1644511149
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1644511149
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1644511149
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1644511149
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_81
timestamp 1644511149
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_93
timestamp 1644511149
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1644511149
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1644511149
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_113
timestamp 1644511149
transform 1 0 11500 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_121
timestamp 1644511149
transform 1 0 12236 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_139
timestamp 1644511149
transform 1 0 13892 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_159
timestamp 1644511149
transform 1 0 15732 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1644511149
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_173
timestamp 1644511149
transform 1 0 17020 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_87_200
timestamp 1644511149
transform 1 0 19504 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_209
timestamp 1644511149
transform 1 0 20332 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_221
timestamp 1644511149
transform 1 0 21436 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_87_225
timestamp 1644511149
transform 1 0 21804 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_231
timestamp 1644511149
transform 1 0 22356 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_253
timestamp 1644511149
transform 1 0 24380 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_261
timestamp 1644511149
transform 1 0 25116 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_269
timestamp 1644511149
transform 1 0 25852 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_87_274
timestamp 1644511149
transform 1 0 26312 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_87_281
timestamp 1644511149
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_293
timestamp 1644511149
transform 1 0 28060 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_87_302
timestamp 1644511149
transform 1 0 28888 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_312
timestamp 1644511149
transform 1 0 29808 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_332
timestamp 1644511149
transform 1 0 31648 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_353
timestamp 1644511149
transform 1 0 33580 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_359
timestamp 1644511149
transform 1 0 34132 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_367
timestamp 1644511149
transform 1 0 34868 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_377
timestamp 1644511149
transform 1 0 35788 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_87_388
timestamp 1644511149
transform 1 0 36800 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_397
timestamp 1644511149
transform 1 0 37628 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_87_407
timestamp 1644511149
transform 1 0 38548 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_428
timestamp 1644511149
transform 1 0 40480 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_444
timestamp 1644511149
transform 1 0 41952 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_453
timestamp 1644511149
transform 1 0 42780 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_87_465
timestamp 1644511149
transform 1 0 43884 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_471
timestamp 1644511149
transform 1 0 44436 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_480
timestamp 1644511149
transform 1 0 45264 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_486
timestamp 1644511149
transform 1 0 45816 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_494
timestamp 1644511149
transform 1 0 46552 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_502
timestamp 1644511149
transform 1 0 47288 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_505
timestamp 1644511149
transform 1 0 47564 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_514
timestamp 1644511149
transform 1 0 48392 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_523
timestamp 1644511149
transform 1 0 49220 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_531
timestamp 1644511149
transform 1 0 49956 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_538
timestamp 1644511149
transform 1 0 50600 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_544
timestamp 1644511149
transform 1 0 51152 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_548
timestamp 1644511149
transform 1 0 51520 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_555
timestamp 1644511149
transform 1 0 52164 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1644511149
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_561
timestamp 1644511149
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_573
timestamp 1644511149
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_585
timestamp 1644511149
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_597
timestamp 1644511149
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1644511149
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1644511149
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_617
timestamp 1644511149
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_629
timestamp 1644511149
transform 1 0 58972 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_641
timestamp 1644511149
transform 1 0 60076 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_653
timestamp 1644511149
transform 1 0 61180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_665
timestamp 1644511149
transform 1 0 62284 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_671
timestamp 1644511149
transform 1 0 62836 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_673
timestamp 1644511149
transform 1 0 63020 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_685
timestamp 1644511149
transform 1 0 64124 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_697
timestamp 1644511149
transform 1 0 65228 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_709
timestamp 1644511149
transform 1 0 66332 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_721
timestamp 1644511149
transform 1 0 67436 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_727
timestamp 1644511149
transform 1 0 67988 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_729
timestamp 1644511149
transform 1 0 68172 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1644511149
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1644511149
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1644511149
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_29
timestamp 1644511149
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_41
timestamp 1644511149
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_53
timestamp 1644511149
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_65
timestamp 1644511149
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1644511149
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1644511149
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_85
timestamp 1644511149
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_97
timestamp 1644511149
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_109
timestamp 1644511149
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_88_121
timestamp 1644511149
transform 1 0 12236 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_88_127
timestamp 1644511149
transform 1 0 12788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1644511149
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_141
timestamp 1644511149
transform 1 0 14076 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_149
timestamp 1644511149
transform 1 0 14812 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_88_156
timestamp 1644511149
transform 1 0 15456 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_88_168
timestamp 1644511149
transform 1 0 16560 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_174
timestamp 1644511149
transform 1 0 17112 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_186
timestamp 1644511149
transform 1 0 18216 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_194
timestamp 1644511149
transform 1 0 18952 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_213
timestamp 1644511149
transform 1 0 20700 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_227
timestamp 1644511149
transform 1 0 21988 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_239
timestamp 1644511149
transform 1 0 23092 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_243
timestamp 1644511149
transform 1 0 23460 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_248
timestamp 1644511149
transform 1 0 23920 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_274
timestamp 1644511149
transform 1 0 26312 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_88_286
timestamp 1644511149
transform 1 0 27416 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_88_291
timestamp 1644511149
transform 1 0 27876 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_303
timestamp 1644511149
transform 1 0 28980 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1644511149
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_309
timestamp 1644511149
transform 1 0 29532 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_323
timestamp 1644511149
transform 1 0 30820 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_335
timestamp 1644511149
transform 1 0 31924 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_88_343
timestamp 1644511149
transform 1 0 32660 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_88_353
timestamp 1644511149
transform 1 0 33580 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_361
timestamp 1644511149
transform 1 0 34316 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_365
timestamp 1644511149
transform 1 0 34684 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_375
timestamp 1644511149
transform 1 0 35604 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_379
timestamp 1644511149
transform 1 0 35972 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_390
timestamp 1644511149
transform 1 0 36984 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_394
timestamp 1644511149
transform 1 0 37352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_401
timestamp 1644511149
transform 1 0 37996 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_405
timestamp 1644511149
transform 1 0 38364 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_88_410
timestamp 1644511149
transform 1 0 38824 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_418
timestamp 1644511149
transform 1 0 39560 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_421
timestamp 1644511149
transform 1 0 39836 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_426
timestamp 1644511149
transform 1 0 40296 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_440
timestamp 1644511149
transform 1 0 41584 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_452
timestamp 1644511149
transform 1 0 42688 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_464
timestamp 1644511149
transform 1 0 43792 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_477
timestamp 1644511149
transform 1 0 44988 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_483
timestamp 1644511149
transform 1 0 45540 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_491
timestamp 1644511149
transform 1 0 46276 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_88_506
timestamp 1644511149
transform 1 0 47656 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_520
timestamp 1644511149
transform 1 0 48944 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_88_533
timestamp 1644511149
transform 1 0 50140 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_88_540
timestamp 1644511149
transform 1 0 50784 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_564
timestamp 1644511149
transform 1 0 52992 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_576
timestamp 1644511149
transform 1 0 54096 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_589
timestamp 1644511149
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_601
timestamp 1644511149
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_613
timestamp 1644511149
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_625
timestamp 1644511149
transform 1 0 58604 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_637
timestamp 1644511149
transform 1 0 59708 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_643
timestamp 1644511149
transform 1 0 60260 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_645
timestamp 1644511149
transform 1 0 60444 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_657
timestamp 1644511149
transform 1 0 61548 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_669
timestamp 1644511149
transform 1 0 62652 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_681
timestamp 1644511149
transform 1 0 63756 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_693
timestamp 1644511149
transform 1 0 64860 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_699
timestamp 1644511149
transform 1 0 65412 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_701
timestamp 1644511149
transform 1 0 65596 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_713
timestamp 1644511149
transform 1 0 66700 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_725
timestamp 1644511149
transform 1 0 67804 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_3
timestamp 1644511149
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_15
timestamp 1644511149
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_27
timestamp 1644511149
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_39
timestamp 1644511149
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1644511149
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1644511149
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1644511149
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1644511149
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_81
timestamp 1644511149
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_93
timestamp 1644511149
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1644511149
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1644511149
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_113
timestamp 1644511149
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_125
timestamp 1644511149
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_137
timestamp 1644511149
transform 1 0 13708 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_143
timestamp 1644511149
transform 1 0 14260 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_150
timestamp 1644511149
transform 1 0 14904 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_162
timestamp 1644511149
transform 1 0 16008 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_89_173
timestamp 1644511149
transform 1 0 17020 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_180
timestamp 1644511149
transform 1 0 17664 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_192
timestamp 1644511149
transform 1 0 18768 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_203
timestamp 1644511149
transform 1 0 19780 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_219
timestamp 1644511149
transform 1 0 21252 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1644511149
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_225
timestamp 1644511149
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_237
timestamp 1644511149
transform 1 0 22908 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_89_249
timestamp 1644511149
transform 1 0 24012 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_257
timestamp 1644511149
transform 1 0 24748 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_89_268
timestamp 1644511149
transform 1 0 25760 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_276
timestamp 1644511149
transform 1 0 26496 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_297
timestamp 1644511149
transform 1 0 28428 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_309
timestamp 1644511149
transform 1 0 29532 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_89_316
timestamp 1644511149
transform 1 0 30176 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_322
timestamp 1644511149
transform 1 0 30728 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_327
timestamp 1644511149
transform 1 0 31188 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1644511149
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_337
timestamp 1644511149
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_349
timestamp 1644511149
transform 1 0 33212 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_357
timestamp 1644511149
transform 1 0 33948 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_89_363
timestamp 1644511149
transform 1 0 34500 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_371
timestamp 1644511149
transform 1 0 35236 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_379
timestamp 1644511149
transform 1 0 35972 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_387
timestamp 1644511149
transform 1 0 36708 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1644511149
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_393
timestamp 1644511149
transform 1 0 37260 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_403
timestamp 1644511149
transform 1 0 38180 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_410
timestamp 1644511149
transform 1 0 38824 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_416
timestamp 1644511149
transform 1 0 39376 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_421
timestamp 1644511149
transform 1 0 39836 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1644511149
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1644511149
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_449
timestamp 1644511149
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_468
timestamp 1644511149
transform 1 0 44160 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_474
timestamp 1644511149
transform 1 0 44712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_485
timestamp 1644511149
transform 1 0 45724 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_496
timestamp 1644511149
transform 1 0 46736 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_89_509
timestamp 1644511149
transform 1 0 47932 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_89_522
timestamp 1644511149
transform 1 0 49128 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_89_540
timestamp 1644511149
transform 1 0 50784 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_544
timestamp 1644511149
transform 1 0 51152 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_550
timestamp 1644511149
transform 1 0 51704 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_558
timestamp 1644511149
transform 1 0 52440 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_564
timestamp 1644511149
transform 1 0 52992 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_576
timestamp 1644511149
transform 1 0 54096 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_588
timestamp 1644511149
transform 1 0 55200 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_600
timestamp 1644511149
transform 1 0 56304 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_612
timestamp 1644511149
transform 1 0 57408 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_617
timestamp 1644511149
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_629
timestamp 1644511149
transform 1 0 58972 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_641
timestamp 1644511149
transform 1 0 60076 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_653
timestamp 1644511149
transform 1 0 61180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_665
timestamp 1644511149
transform 1 0 62284 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_671
timestamp 1644511149
transform 1 0 62836 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_673
timestamp 1644511149
transform 1 0 63020 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_685
timestamp 1644511149
transform 1 0 64124 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_697
timestamp 1644511149
transform 1 0 65228 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_712
timestamp 1644511149
transform 1 0 66608 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_724
timestamp 1644511149
transform 1 0 67712 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_729
timestamp 1644511149
transform 1 0 68172 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1644511149
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1644511149
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1644511149
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1644511149
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_41
timestamp 1644511149
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_53
timestamp 1644511149
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_65
timestamp 1644511149
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1644511149
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1644511149
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_85
timestamp 1644511149
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_97
timestamp 1644511149
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_109
timestamp 1644511149
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_121
timestamp 1644511149
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1644511149
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1644511149
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_141
timestamp 1644511149
transform 1 0 14076 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_146
timestamp 1644511149
transform 1 0 14536 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_150
timestamp 1644511149
transform 1 0 14904 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_154
timestamp 1644511149
transform 1 0 15272 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_163
timestamp 1644511149
transform 1 0 16100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_169
timestamp 1644511149
transform 1 0 16652 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_186
timestamp 1644511149
transform 1 0 18216 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_194
timestamp 1644511149
transform 1 0 18952 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_197
timestamp 1644511149
transform 1 0 19228 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_201
timestamp 1644511149
transform 1 0 19596 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_205
timestamp 1644511149
transform 1 0 19964 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_209
timestamp 1644511149
transform 1 0 20332 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_214
timestamp 1644511149
transform 1 0 20792 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_232
timestamp 1644511149
transform 1 0 22448 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_248
timestamp 1644511149
transform 1 0 23920 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_253
timestamp 1644511149
transform 1 0 24380 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_257
timestamp 1644511149
transform 1 0 24748 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_274
timestamp 1644511149
transform 1 0 26312 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_281
timestamp 1644511149
transform 1 0 26956 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_90_289
timestamp 1644511149
transform 1 0 27692 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_90_302
timestamp 1644511149
transform 1 0 28888 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_90_330
timestamp 1644511149
transform 1 0 31464 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_342
timestamp 1644511149
transform 1 0 32568 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_360
timestamp 1644511149
transform 1 0 34224 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_368
timestamp 1644511149
transform 1 0 34960 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_372
timestamp 1644511149
transform 1 0 35328 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_380
timestamp 1644511149
transform 1 0 36064 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_388
timestamp 1644511149
transform 1 0 36800 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_402
timestamp 1644511149
transform 1 0 38088 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_412
timestamp 1644511149
transform 1 0 39008 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_90_437
timestamp 1644511149
transform 1 0 41308 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_445
timestamp 1644511149
transform 1 0 42044 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_457
timestamp 1644511149
transform 1 0 43148 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_468
timestamp 1644511149
transform 1 0 44160 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_90_480
timestamp 1644511149
transform 1 0 45264 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_491
timestamp 1644511149
transform 1 0 46276 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_503
timestamp 1644511149
transform 1 0 47380 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_515
timestamp 1644511149
transform 1 0 48484 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_90_528
timestamp 1644511149
transform 1 0 49680 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_533
timestamp 1644511149
transform 1 0 50140 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_539
timestamp 1644511149
transform 1 0 50692 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_546
timestamp 1644511149
transform 1 0 51336 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_558
timestamp 1644511149
transform 1 0 52440 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_570
timestamp 1644511149
transform 1 0 53544 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_582
timestamp 1644511149
transform 1 0 54648 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_90_589
timestamp 1644511149
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_601
timestamp 1644511149
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_613
timestamp 1644511149
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_625
timestamp 1644511149
transform 1 0 58604 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_637
timestamp 1644511149
transform 1 0 59708 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_643
timestamp 1644511149
transform 1 0 60260 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_645
timestamp 1644511149
transform 1 0 60444 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_657
timestamp 1644511149
transform 1 0 61548 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_669
timestamp 1644511149
transform 1 0 62652 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_681
timestamp 1644511149
transform 1 0 63756 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_693
timestamp 1644511149
transform 1 0 64860 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_699
timestamp 1644511149
transform 1 0 65412 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_701
timestamp 1644511149
transform 1 0 65596 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_707
timestamp 1644511149
transform 1 0 66148 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_729
timestamp 1644511149
transform 1 0 68172 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_91_3
timestamp 1644511149
transform 1 0 1380 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_91_12
timestamp 1644511149
transform 1 0 2208 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_24
timestamp 1644511149
transform 1 0 3312 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_36
timestamp 1644511149
transform 1 0 4416 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_48
timestamp 1644511149
transform 1 0 5520 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1644511149
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1644511149
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_81
timestamp 1644511149
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_93
timestamp 1644511149
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1644511149
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1644511149
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_113
timestamp 1644511149
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_125
timestamp 1644511149
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_137
timestamp 1644511149
transform 1 0 13708 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_143
timestamp 1644511149
transform 1 0 14260 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_160
timestamp 1644511149
transform 1 0 15824 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_91_169
timestamp 1644511149
transform 1 0 16652 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_91_198
timestamp 1644511149
transform 1 0 19320 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_91_207
timestamp 1644511149
transform 1 0 20148 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_213
timestamp 1644511149
transform 1 0 20700 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_91_218
timestamp 1644511149
transform 1 0 21160 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_91_241
timestamp 1644511149
transform 1 0 23276 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_253
timestamp 1644511149
transform 1 0 24380 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_91_271
timestamp 1644511149
transform 1 0 26036 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1644511149
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_281
timestamp 1644511149
transform 1 0 26956 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_289
timestamp 1644511149
transform 1 0 27692 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_91_297
timestamp 1644511149
transform 1 0 28428 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_305
timestamp 1644511149
transform 1 0 29164 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_317
timestamp 1644511149
transform 1 0 30268 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_331
timestamp 1644511149
transform 1 0 31556 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1644511149
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_342
timestamp 1644511149
transform 1 0 32568 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_354
timestamp 1644511149
transform 1 0 33672 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_366
timestamp 1644511149
transform 1 0 34776 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_375
timestamp 1644511149
transform 1 0 35604 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_387
timestamp 1644511149
transform 1 0 36708 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1644511149
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_91_393
timestamp 1644511149
transform 1 0 37260 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_91_416
timestamp 1644511149
transform 1 0 39376 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_428
timestamp 1644511149
transform 1 0 40480 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_91_444
timestamp 1644511149
transform 1 0 41952 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_455
timestamp 1644511149
transform 1 0 42964 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_468
timestamp 1644511149
transform 1 0 44160 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_480
timestamp 1644511149
transform 1 0 45264 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_91_494
timestamp 1644511149
transform 1 0 46552 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_502
timestamp 1644511149
transform 1 0 47288 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_91_521
timestamp 1644511149
transform 1 0 49036 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_545
timestamp 1644511149
transform 1 0 51244 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_557
timestamp 1644511149
transform 1 0 52348 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_561
timestamp 1644511149
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_573
timestamp 1644511149
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_585
timestamp 1644511149
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_597
timestamp 1644511149
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1644511149
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1644511149
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_617
timestamp 1644511149
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_629
timestamp 1644511149
transform 1 0 58972 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_641
timestamp 1644511149
transform 1 0 60076 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_653
timestamp 1644511149
transform 1 0 61180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_665
timestamp 1644511149
transform 1 0 62284 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_671
timestamp 1644511149
transform 1 0 62836 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_673
timestamp 1644511149
transform 1 0 63020 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_685
timestamp 1644511149
transform 1 0 64124 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_697
timestamp 1644511149
transform 1 0 65228 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_709
timestamp 1644511149
transform 1 0 66332 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_717
timestamp 1644511149
transform 1 0 67068 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_91_721
timestamp 1644511149
transform 1 0 67436 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_727
timestamp 1644511149
transform 1 0 67988 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_729
timestamp 1644511149
transform 1 0 68172 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_24
timestamp 1644511149
transform 1 0 3312 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_29
timestamp 1644511149
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_41
timestamp 1644511149
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_53
timestamp 1644511149
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_65
timestamp 1644511149
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1644511149
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1644511149
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_85
timestamp 1644511149
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_97
timestamp 1644511149
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_109
timestamp 1644511149
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_121
timestamp 1644511149
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1644511149
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1644511149
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_144
timestamp 1644511149
transform 1 0 14352 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_156
timestamp 1644511149
transform 1 0 15456 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_160
timestamp 1644511149
transform 1 0 15824 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_165
timestamp 1644511149
transform 1 0 16284 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_179
timestamp 1644511149
transform 1 0 17572 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_188
timestamp 1644511149
transform 1 0 18400 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_197
timestamp 1644511149
transform 1 0 19228 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_214
timestamp 1644511149
transform 1 0 20792 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_92_228
timestamp 1644511149
transform 1 0 22080 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_248
timestamp 1644511149
transform 1 0 23920 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_253
timestamp 1644511149
transform 1 0 24380 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_258
timestamp 1644511149
transform 1 0 24840 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_265
timestamp 1644511149
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_277
timestamp 1644511149
transform 1 0 26588 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_295
timestamp 1644511149
transform 1 0 28244 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_304
timestamp 1644511149
transform 1 0 29072 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_313
timestamp 1644511149
transform 1 0 29900 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_317
timestamp 1644511149
transform 1 0 30268 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_322
timestamp 1644511149
transform 1 0 30728 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_342
timestamp 1644511149
transform 1 0 32568 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_350
timestamp 1644511149
transform 1 0 33304 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_92_356
timestamp 1644511149
transform 1 0 33856 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_92_365
timestamp 1644511149
transform 1 0 34684 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_376
timestamp 1644511149
transform 1 0 35696 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_388
timestamp 1644511149
transform 1 0 36800 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_400
timestamp 1644511149
transform 1 0 37904 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_412
timestamp 1644511149
transform 1 0 39008 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_421
timestamp 1644511149
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_433
timestamp 1644511149
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_445
timestamp 1644511149
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_457
timestamp 1644511149
transform 1 0 43148 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_92_472
timestamp 1644511149
transform 1 0 44528 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_477
timestamp 1644511149
transform 1 0 44988 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_485
timestamp 1644511149
transform 1 0 45724 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_496
timestamp 1644511149
transform 1 0 46736 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_504
timestamp 1644511149
transform 1 0 47472 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_509
timestamp 1644511149
transform 1 0 47932 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_521
timestamp 1644511149
transform 1 0 49036 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_529
timestamp 1644511149
transform 1 0 49772 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_537
timestamp 1644511149
transform 1 0 50508 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_549
timestamp 1644511149
transform 1 0 51612 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_561
timestamp 1644511149
transform 1 0 52716 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_573
timestamp 1644511149
transform 1 0 53820 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_585
timestamp 1644511149
transform 1 0 54924 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_589
timestamp 1644511149
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_601
timestamp 1644511149
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_613
timestamp 1644511149
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_625
timestamp 1644511149
transform 1 0 58604 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_637
timestamp 1644511149
transform 1 0 59708 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_643
timestamp 1644511149
transform 1 0 60260 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_645
timestamp 1644511149
transform 1 0 60444 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_657
timestamp 1644511149
transform 1 0 61548 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_669
timestamp 1644511149
transform 1 0 62652 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_681
timestamp 1644511149
transform 1 0 63756 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_693
timestamp 1644511149
transform 1 0 64860 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_699
timestamp 1644511149
transform 1 0 65412 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_701
timestamp 1644511149
transform 1 0 65596 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_713
timestamp 1644511149
transform 1 0 66700 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_725
timestamp 1644511149
transform 1 0 67804 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1644511149
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_8
timestamp 1644511149
transform 1 0 1840 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_12
timestamp 1644511149
transform 1 0 2208 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_16
timestamp 1644511149
transform 1 0 2576 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_28
timestamp 1644511149
transform 1 0 3680 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_40
timestamp 1644511149
transform 1 0 4784 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_52
timestamp 1644511149
transform 1 0 5888 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_57
timestamp 1644511149
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_69
timestamp 1644511149
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_81
timestamp 1644511149
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_93
timestamp 1644511149
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1644511149
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1644511149
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_113
timestamp 1644511149
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_125
timestamp 1644511149
transform 1 0 12604 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_133
timestamp 1644511149
transform 1 0 13340 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_151
timestamp 1644511149
transform 1 0 14996 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1644511149
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1644511149
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_172
timestamp 1644511149
transform 1 0 16928 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_184
timestamp 1644511149
transform 1 0 18032 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_196
timestamp 1644511149
transform 1 0 19136 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_202
timestamp 1644511149
transform 1 0 19688 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_218
timestamp 1644511149
transform 1 0 21160 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_93_225
timestamp 1644511149
transform 1 0 21804 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_93_241
timestamp 1644511149
transform 1 0 23276 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_249
timestamp 1644511149
transform 1 0 24012 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_258
timestamp 1644511149
transform 1 0 24840 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_262
timestamp 1644511149
transform 1 0 25208 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_268
timestamp 1644511149
transform 1 0 25760 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_281
timestamp 1644511149
transform 1 0 26956 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_285
timestamp 1644511149
transform 1 0 27324 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_289
timestamp 1644511149
transform 1 0 27692 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_93_314
timestamp 1644511149
transform 1 0 29992 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_322
timestamp 1644511149
transform 1 0 30728 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_327
timestamp 1644511149
transform 1 0 31188 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1644511149
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_337
timestamp 1644511149
transform 1 0 32108 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_345
timestamp 1644511149
transform 1 0 32844 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_93_364
timestamp 1644511149
transform 1 0 34592 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_93_381
timestamp 1644511149
transform 1 0 36156 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_389
timestamp 1644511149
transform 1 0 36892 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_399
timestamp 1644511149
transform 1 0 37812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_411
timestamp 1644511149
transform 1 0 38916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_433
timestamp 1644511149
transform 1 0 40940 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_444
timestamp 1644511149
transform 1 0 41952 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_453
timestamp 1644511149
transform 1 0 42780 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_457
timestamp 1644511149
transform 1 0 43148 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_462
timestamp 1644511149
transform 1 0 43608 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_474
timestamp 1644511149
transform 1 0 44712 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_485
timestamp 1644511149
transform 1 0 45724 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_93_495
timestamp 1644511149
transform 1 0 46644 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1644511149
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_513
timestamp 1644511149
transform 1 0 48300 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_525
timestamp 1644511149
transform 1 0 49404 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_529
timestamp 1644511149
transform 1 0 49772 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_535
timestamp 1644511149
transform 1 0 50324 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_543
timestamp 1644511149
transform 1 0 51060 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_555
timestamp 1644511149
transform 1 0 52164 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1644511149
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_561
timestamp 1644511149
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_573
timestamp 1644511149
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_585
timestamp 1644511149
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_597
timestamp 1644511149
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1644511149
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1644511149
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_617
timestamp 1644511149
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_629
timestamp 1644511149
transform 1 0 58972 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_641
timestamp 1644511149
transform 1 0 60076 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_653
timestamp 1644511149
transform 1 0 61180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_665
timestamp 1644511149
transform 1 0 62284 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_671
timestamp 1644511149
transform 1 0 62836 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_673
timestamp 1644511149
transform 1 0 63020 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_685
timestamp 1644511149
transform 1 0 64124 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_697
timestamp 1644511149
transform 1 0 65228 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_709
timestamp 1644511149
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_721
timestamp 1644511149
transform 1 0 67436 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_727
timestamp 1644511149
transform 1 0 67988 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_729
timestamp 1644511149
transform 1 0 68172 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_24
timestamp 1644511149
transform 1 0 3312 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1644511149
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1644511149
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_56
timestamp 1644511149
transform 1 0 6256 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_68
timestamp 1644511149
transform 1 0 7360 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_80
timestamp 1644511149
transform 1 0 8464 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_85
timestamp 1644511149
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_97
timestamp 1644511149
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_109
timestamp 1644511149
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_121
timestamp 1644511149
transform 1 0 12236 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_129
timestamp 1644511149
transform 1 0 12972 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_136
timestamp 1644511149
transform 1 0 13616 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_141
timestamp 1644511149
transform 1 0 14076 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_150
timestamp 1644511149
transform 1 0 14904 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_156
timestamp 1644511149
transform 1 0 15456 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_173
timestamp 1644511149
transform 1 0 17020 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_181
timestamp 1644511149
transform 1 0 17756 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_187
timestamp 1644511149
transform 1 0 18308 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_192
timestamp 1644511149
transform 1 0 18768 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_197
timestamp 1644511149
transform 1 0 19228 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_94_208
timestamp 1644511149
transform 1 0 20240 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_94_220
timestamp 1644511149
transform 1 0 21344 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_228
timestamp 1644511149
transform 1 0 22080 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_242
timestamp 1644511149
transform 1 0 23368 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1644511149
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_253
timestamp 1644511149
transform 1 0 24380 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_257
timestamp 1644511149
transform 1 0 24748 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_274
timestamp 1644511149
transform 1 0 26312 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_280
timestamp 1644511149
transform 1 0 26864 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_284
timestamp 1644511149
transform 1 0 27232 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_293
timestamp 1644511149
transform 1 0 28060 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_305
timestamp 1644511149
transform 1 0 29164 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_94_309
timestamp 1644511149
transform 1 0 29532 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_317
timestamp 1644511149
transform 1 0 30268 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_324
timestamp 1644511149
transform 1 0 30912 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_330
timestamp 1644511149
transform 1 0 31464 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_341
timestamp 1644511149
transform 1 0 32476 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_353
timestamp 1644511149
transform 1 0 33580 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_361
timestamp 1644511149
transform 1 0 34316 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_365
timestamp 1644511149
transform 1 0 34684 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_375
timestamp 1644511149
transform 1 0 35604 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_383
timestamp 1644511149
transform 1 0 36340 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_94_401
timestamp 1644511149
transform 1 0 37996 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_409
timestamp 1644511149
transform 1 0 38732 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_416
timestamp 1644511149
transform 1 0 39376 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_421
timestamp 1644511149
transform 1 0 39836 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_431
timestamp 1644511149
transform 1 0 40756 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_94_455
timestamp 1644511149
transform 1 0 42964 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_461
timestamp 1644511149
transform 1 0 43516 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_465
timestamp 1644511149
transform 1 0 43884 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_473
timestamp 1644511149
transform 1 0 44620 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_94_477
timestamp 1644511149
transform 1 0 44988 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_482
timestamp 1644511149
transform 1 0 45448 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_493
timestamp 1644511149
transform 1 0 46460 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_505
timestamp 1644511149
transform 1 0 47564 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_94_521
timestamp 1644511149
transform 1 0 49036 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_529
timestamp 1644511149
transform 1 0 49772 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_533
timestamp 1644511149
transform 1 0 50140 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_553
timestamp 1644511149
transform 1 0 51980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_565
timestamp 1644511149
transform 1 0 53084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_577
timestamp 1644511149
transform 1 0 54188 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_585
timestamp 1644511149
transform 1 0 54924 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_589
timestamp 1644511149
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_601
timestamp 1644511149
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_613
timestamp 1644511149
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_625
timestamp 1644511149
transform 1 0 58604 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_637
timestamp 1644511149
transform 1 0 59708 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_643
timestamp 1644511149
transform 1 0 60260 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_645
timestamp 1644511149
transform 1 0 60444 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_657
timestamp 1644511149
transform 1 0 61548 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_669
timestamp 1644511149
transform 1 0 62652 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_681
timestamp 1644511149
transform 1 0 63756 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_693
timestamp 1644511149
transform 1 0 64860 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_699
timestamp 1644511149
transform 1 0 65412 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_701
timestamp 1644511149
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_713
timestamp 1644511149
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_725
timestamp 1644511149
transform 1 0 67804 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_95_3
timestamp 1644511149
transform 1 0 1380 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_10
timestamp 1644511149
transform 1 0 2024 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_22
timestamp 1644511149
transform 1 0 3128 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_34
timestamp 1644511149
transform 1 0 4232 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_46
timestamp 1644511149
transform 1 0 5336 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1644511149
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_95_78
timestamp 1644511149
transform 1 0 8280 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_90
timestamp 1644511149
transform 1 0 9384 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_102
timestamp 1644511149
transform 1 0 10488 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1644511149
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_95_113
timestamp 1644511149
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_125
timestamp 1644511149
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_137
timestamp 1644511149
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_149
timestamp 1644511149
transform 1 0 14812 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_157
timestamp 1644511149
transform 1 0 15548 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_164
timestamp 1644511149
transform 1 0 16192 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_169
timestamp 1644511149
transform 1 0 16652 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_175
timestamp 1644511149
transform 1 0 17204 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_197
timestamp 1644511149
transform 1 0 19228 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1644511149
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1644511149
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_231
timestamp 1644511149
transform 1 0 22356 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_239
timestamp 1644511149
transform 1 0 23092 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_256
timestamp 1644511149
transform 1 0 24656 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_264
timestamp 1644511149
transform 1 0 25392 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_95_276
timestamp 1644511149
transform 1 0 26496 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_297
timestamp 1644511149
transform 1 0 28428 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_309
timestamp 1644511149
transform 1 0 29532 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_328
timestamp 1644511149
transform 1 0 31280 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_354
timestamp 1644511149
transform 1 0 33672 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_366
timestamp 1644511149
transform 1 0 34776 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_378
timestamp 1644511149
transform 1 0 35880 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_390
timestamp 1644511149
transform 1 0 36984 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_393
timestamp 1644511149
transform 1 0 37260 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_412
timestamp 1644511149
transform 1 0 39008 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_420
timestamp 1644511149
transform 1 0 39744 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_427
timestamp 1644511149
transform 1 0 40388 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_434
timestamp 1644511149
transform 1 0 41032 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1644511149
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1644511149
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_449
timestamp 1644511149
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_95_461
timestamp 1644511149
transform 1 0 43516 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_478
timestamp 1644511149
transform 1 0 45080 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_95_490
timestamp 1644511149
transform 1 0 46184 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_502
timestamp 1644511149
transform 1 0 47288 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_509
timestamp 1644511149
transform 1 0 47932 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_515
timestamp 1644511149
transform 1 0 48484 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_521
timestamp 1644511149
transform 1 0 49036 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_529
timestamp 1644511149
transform 1 0 49772 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_535
timestamp 1644511149
transform 1 0 50324 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_542
timestamp 1644511149
transform 1 0 50968 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_554
timestamp 1644511149
transform 1 0 52072 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_95_561
timestamp 1644511149
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_573
timestamp 1644511149
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_585
timestamp 1644511149
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_597
timestamp 1644511149
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1644511149
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1644511149
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_617
timestamp 1644511149
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_629
timestamp 1644511149
transform 1 0 58972 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_641
timestamp 1644511149
transform 1 0 60076 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_653
timestamp 1644511149
transform 1 0 61180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_665
timestamp 1644511149
transform 1 0 62284 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_671
timestamp 1644511149
transform 1 0 62836 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_673
timestamp 1644511149
transform 1 0 63020 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_685
timestamp 1644511149
transform 1 0 64124 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_697
timestamp 1644511149
transform 1 0 65228 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_709
timestamp 1644511149
transform 1 0 66332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_721
timestamp 1644511149
transform 1 0 67436 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_727
timestamp 1644511149
transform 1 0 67988 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_729
timestamp 1644511149
transform 1 0 68172 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_3
timestamp 1644511149
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1644511149
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1644511149
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1644511149
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_41
timestamp 1644511149
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_53
timestamp 1644511149
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_65
timestamp 1644511149
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1644511149
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1644511149
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_85
timestamp 1644511149
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_97
timestamp 1644511149
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_109
timestamp 1644511149
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_121
timestamp 1644511149
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1644511149
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1644511149
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_141
timestamp 1644511149
transform 1 0 14076 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_149
timestamp 1644511149
transform 1 0 14812 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_155
timestamp 1644511149
transform 1 0 15364 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_167
timestamp 1644511149
transform 1 0 16468 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_179
timestamp 1644511149
transform 1 0 17572 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_183
timestamp 1644511149
transform 1 0 17940 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1644511149
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_197
timestamp 1644511149
transform 1 0 19228 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_203
timestamp 1644511149
transform 1 0 19780 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_210
timestamp 1644511149
transform 1 0 20424 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_220
timestamp 1644511149
transform 1 0 21344 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_232
timestamp 1644511149
transform 1 0 22448 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_236
timestamp 1644511149
transform 1 0 22816 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1644511149
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1644511149
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_253
timestamp 1644511149
transform 1 0 24380 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_261
timestamp 1644511149
transform 1 0 25116 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_265
timestamp 1644511149
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_277
timestamp 1644511149
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_289
timestamp 1644511149
transform 1 0 27692 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_96_297
timestamp 1644511149
transform 1 0 28428 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_304
timestamp 1644511149
transform 1 0 29072 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_309
timestamp 1644511149
transform 1 0 29532 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_317
timestamp 1644511149
transform 1 0 30268 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_335
timestamp 1644511149
transform 1 0 31924 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_343
timestamp 1644511149
transform 1 0 32660 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_355
timestamp 1644511149
transform 1 0 33764 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1644511149
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_371
timestamp 1644511149
transform 1 0 35236 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_379
timestamp 1644511149
transform 1 0 35972 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_391
timestamp 1644511149
transform 1 0 37076 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_403
timestamp 1644511149
transform 1 0 38180 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_410
timestamp 1644511149
transform 1 0 38824 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_418
timestamp 1644511149
transform 1 0 39560 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_96_421
timestamp 1644511149
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_433
timestamp 1644511149
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_445
timestamp 1644511149
transform 1 0 42044 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_453
timestamp 1644511149
transform 1 0 42780 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_458
timestamp 1644511149
transform 1 0 43240 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_466
timestamp 1644511149
transform 1 0 43976 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_471
timestamp 1644511149
transform 1 0 44436 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1644511149
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_481
timestamp 1644511149
transform 1 0 45356 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_501
timestamp 1644511149
transform 1 0 47196 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_505
timestamp 1644511149
transform 1 0 47564 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_522
timestamp 1644511149
transform 1 0 49128 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_530
timestamp 1644511149
transform 1 0 49864 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_96_533
timestamp 1644511149
transform 1 0 50140 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_552
timestamp 1644511149
transform 1 0 51888 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_564
timestamp 1644511149
transform 1 0 52992 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_576
timestamp 1644511149
transform 1 0 54096 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_589
timestamp 1644511149
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_601
timestamp 1644511149
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_613
timestamp 1644511149
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_625
timestamp 1644511149
transform 1 0 58604 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_637
timestamp 1644511149
transform 1 0 59708 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_643
timestamp 1644511149
transform 1 0 60260 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_645
timestamp 1644511149
transform 1 0 60444 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_657
timestamp 1644511149
transform 1 0 61548 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_669
timestamp 1644511149
transform 1 0 62652 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_681
timestamp 1644511149
transform 1 0 63756 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_693
timestamp 1644511149
transform 1 0 64860 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_699
timestamp 1644511149
transform 1 0 65412 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_701
timestamp 1644511149
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_713
timestamp 1644511149
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_725
timestamp 1644511149
transform 1 0 67804 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1644511149
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1644511149
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1644511149
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1644511149
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1644511149
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1644511149
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1644511149
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1644511149
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_81
timestamp 1644511149
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_93
timestamp 1644511149
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1644511149
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1644511149
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_113
timestamp 1644511149
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_125
timestamp 1644511149
transform 1 0 12604 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_133
timestamp 1644511149
transform 1 0 13340 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_138
timestamp 1644511149
transform 1 0 13800 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_158
timestamp 1644511149
transform 1 0 15640 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_166
timestamp 1644511149
transform 1 0 16376 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_97_169
timestamp 1644511149
transform 1 0 16652 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_188
timestamp 1644511149
transform 1 0 18400 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_197
timestamp 1644511149
transform 1 0 19228 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_209
timestamp 1644511149
transform 1 0 20332 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_221
timestamp 1644511149
transform 1 0 21436 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_225
timestamp 1644511149
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_237
timestamp 1644511149
transform 1 0 22908 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_246
timestamp 1644511149
transform 1 0 23736 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_258
timestamp 1644511149
transform 1 0 24840 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_265
timestamp 1644511149
transform 1 0 25484 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_277
timestamp 1644511149
transform 1 0 26588 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_97_281
timestamp 1644511149
transform 1 0 26956 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_97_291
timestamp 1644511149
transform 1 0 27876 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_297
timestamp 1644511149
transform 1 0 28428 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_301
timestamp 1644511149
transform 1 0 28796 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_313
timestamp 1644511149
transform 1 0 29900 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_325
timestamp 1644511149
transform 1 0 31004 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_332
timestamp 1644511149
transform 1 0 31648 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_337
timestamp 1644511149
transform 1 0 32108 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_341
timestamp 1644511149
transform 1 0 32476 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_345
timestamp 1644511149
transform 1 0 32844 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_97_369
timestamp 1644511149
transform 1 0 35052 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_97_380
timestamp 1644511149
transform 1 0 36064 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_384
timestamp 1644511149
transform 1 0 36432 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_388
timestamp 1644511149
transform 1 0 36800 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_393
timestamp 1644511149
transform 1 0 37260 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_97_403
timestamp 1644511149
transform 1 0 38180 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_97_415
timestamp 1644511149
transform 1 0 39284 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_427
timestamp 1644511149
transform 1 0 40388 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_434
timestamp 1644511149
transform 1 0 41032 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_446
timestamp 1644511149
transform 1 0 42136 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_97_449
timestamp 1644511149
transform 1 0 42412 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_466
timestamp 1644511149
transform 1 0 43976 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_478
timestamp 1644511149
transform 1 0 45080 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_484
timestamp 1644511149
transform 1 0 45632 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_489
timestamp 1644511149
transform 1 0 46092 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_501
timestamp 1644511149
transform 1 0 47196 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_508
timestamp 1644511149
transform 1 0 47840 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_512
timestamp 1644511149
transform 1 0 48208 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_516
timestamp 1644511149
transform 1 0 48576 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_528
timestamp 1644511149
transform 1 0 49680 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_534
timestamp 1644511149
transform 1 0 50232 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_539
timestamp 1644511149
transform 1 0 50692 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_546
timestamp 1644511149
transform 1 0 51336 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_558
timestamp 1644511149
transform 1 0 52440 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_561
timestamp 1644511149
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_573
timestamp 1644511149
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_585
timestamp 1644511149
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_597
timestamp 1644511149
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1644511149
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1644511149
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_617
timestamp 1644511149
transform 1 0 57868 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_629
timestamp 1644511149
transform 1 0 58972 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_641
timestamp 1644511149
transform 1 0 60076 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_653
timestamp 1644511149
transform 1 0 61180 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_665
timestamp 1644511149
transform 1 0 62284 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_671
timestamp 1644511149
transform 1 0 62836 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_673
timestamp 1644511149
transform 1 0 63020 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_685
timestamp 1644511149
transform 1 0 64124 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_697
timestamp 1644511149
transform 1 0 65228 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_709
timestamp 1644511149
transform 1 0 66332 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_721
timestamp 1644511149
transform 1 0 67436 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_727
timestamp 1644511149
transform 1 0 67988 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_729
timestamp 1644511149
transform 1 0 68172 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1644511149
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1644511149
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1644511149
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_29
timestamp 1644511149
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_41
timestamp 1644511149
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_53
timestamp 1644511149
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_65
timestamp 1644511149
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1644511149
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1644511149
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_85
timestamp 1644511149
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_97
timestamp 1644511149
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_109
timestamp 1644511149
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_121
timestamp 1644511149
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1644511149
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1644511149
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_141
timestamp 1644511149
transform 1 0 14076 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_98_150
timestamp 1644511149
transform 1 0 14904 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_158
timestamp 1644511149
transform 1 0 15640 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_164
timestamp 1644511149
transform 1 0 16192 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_172
timestamp 1644511149
transform 1 0 16928 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_184
timestamp 1644511149
transform 1 0 18032 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_197
timestamp 1644511149
transform 1 0 19228 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_203
timestamp 1644511149
transform 1 0 19780 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_209
timestamp 1644511149
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_221
timestamp 1644511149
transform 1 0 21436 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_241
timestamp 1644511149
transform 1 0 23276 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_249
timestamp 1644511149
transform 1 0 24012 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_98_253
timestamp 1644511149
transform 1 0 24380 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_270
timestamp 1644511149
transform 1 0 25944 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_98_279
timestamp 1644511149
transform 1 0 26772 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_288
timestamp 1644511149
transform 1 0 27600 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_296
timestamp 1644511149
transform 1 0 28336 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_302
timestamp 1644511149
transform 1 0 28888 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_309
timestamp 1644511149
transform 1 0 29532 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_314
timestamp 1644511149
transform 1 0 29992 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_323
timestamp 1644511149
transform 1 0 30820 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_331
timestamp 1644511149
transform 1 0 31556 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_98_360
timestamp 1644511149
transform 1 0 34224 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_365
timestamp 1644511149
transform 1 0 34684 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_373
timestamp 1644511149
transform 1 0 35420 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_385
timestamp 1644511149
transform 1 0 36524 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_396
timestamp 1644511149
transform 1 0 37536 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_404
timestamp 1644511149
transform 1 0 38272 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_414
timestamp 1644511149
transform 1 0 39192 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_98_421
timestamp 1644511149
transform 1 0 39836 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_440
timestamp 1644511149
transform 1 0 41584 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_452
timestamp 1644511149
transform 1 0 42688 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_464
timestamp 1644511149
transform 1 0 43792 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_482
timestamp 1644511149
transform 1 0 45448 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_489
timestamp 1644511149
transform 1 0 46092 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_98_499
timestamp 1644511149
transform 1 0 47012 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_98_509
timestamp 1644511149
transform 1 0 47932 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_515
timestamp 1644511149
transform 1 0 48484 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_520
timestamp 1644511149
transform 1 0 48944 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_538
timestamp 1644511149
transform 1 0 50600 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_550
timestamp 1644511149
transform 1 0 51704 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_562
timestamp 1644511149
transform 1 0 52808 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_574
timestamp 1644511149
transform 1 0 53912 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_98_586
timestamp 1644511149
transform 1 0 55016 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_98_589
timestamp 1644511149
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_601
timestamp 1644511149
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_613
timestamp 1644511149
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_625
timestamp 1644511149
transform 1 0 58604 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_637
timestamp 1644511149
transform 1 0 59708 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_643
timestamp 1644511149
transform 1 0 60260 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_645
timestamp 1644511149
transform 1 0 60444 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_657
timestamp 1644511149
transform 1 0 61548 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_669
timestamp 1644511149
transform 1 0 62652 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_681
timestamp 1644511149
transform 1 0 63756 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_693
timestamp 1644511149
transform 1 0 64860 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_699
timestamp 1644511149
transform 1 0 65412 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_701
timestamp 1644511149
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_713
timestamp 1644511149
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_725
timestamp 1644511149
transform 1 0 67804 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_3
timestamp 1644511149
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_15
timestamp 1644511149
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_27
timestamp 1644511149
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_39
timestamp 1644511149
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1644511149
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1644511149
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_57
timestamp 1644511149
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_69
timestamp 1644511149
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_81
timestamp 1644511149
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_93
timestamp 1644511149
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1644511149
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1644511149
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_113
timestamp 1644511149
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_125
timestamp 1644511149
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_137
timestamp 1644511149
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_149
timestamp 1644511149
transform 1 0 14812 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_153
timestamp 1644511149
transform 1 0 15180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_165
timestamp 1644511149
transform 1 0 16284 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_185
timestamp 1644511149
transform 1 0 18124 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_197
timestamp 1644511149
transform 1 0 19228 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_201
timestamp 1644511149
transform 1 0 19596 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_218
timestamp 1644511149
transform 1 0 21160 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_231
timestamp 1644511149
transform 1 0 22356 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_243
timestamp 1644511149
transform 1 0 23460 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_259
timestamp 1644511149
transform 1 0 24932 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_266
timestamp 1644511149
transform 1 0 25576 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_274
timestamp 1644511149
transform 1 0 26312 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_99_281
timestamp 1644511149
transform 1 0 26956 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_299
timestamp 1644511149
transform 1 0 28612 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_324
timestamp 1644511149
transform 1 0 30912 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_337
timestamp 1644511149
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_349
timestamp 1644511149
transform 1 0 33212 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_366
timestamp 1644511149
transform 1 0 34776 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_370
timestamp 1644511149
transform 1 0 35144 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_378
timestamp 1644511149
transform 1 0 35880 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_382
timestamp 1644511149
transform 1 0 36248 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_387
timestamp 1644511149
transform 1 0 36708 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1644511149
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_393
timestamp 1644511149
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_405
timestamp 1644511149
transform 1 0 38364 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_411
timestamp 1644511149
transform 1 0 38916 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_419
timestamp 1644511149
transform 1 0 39652 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_427
timestamp 1644511149
transform 1 0 40388 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_433
timestamp 1644511149
transform 1 0 40940 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_445
timestamp 1644511149
transform 1 0 42044 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_455
timestamp 1644511149
transform 1 0 42964 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_465
timestamp 1644511149
transform 1 0 43884 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_477
timestamp 1644511149
transform 1 0 44988 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_99_495
timestamp 1644511149
transform 1 0 46644 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1644511149
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_505
timestamp 1644511149
transform 1 0 47564 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_99_516
timestamp 1644511149
transform 1 0 48576 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_538
timestamp 1644511149
transform 1 0 50600 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_550
timestamp 1644511149
transform 1 0 51704 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_558
timestamp 1644511149
transform 1 0 52440 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_561
timestamp 1644511149
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_573
timestamp 1644511149
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_585
timestamp 1644511149
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_597
timestamp 1644511149
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1644511149
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1644511149
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_617
timestamp 1644511149
transform 1 0 57868 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_629
timestamp 1644511149
transform 1 0 58972 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_641
timestamp 1644511149
transform 1 0 60076 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_653
timestamp 1644511149
transform 1 0 61180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_665
timestamp 1644511149
transform 1 0 62284 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_671
timestamp 1644511149
transform 1 0 62836 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_673
timestamp 1644511149
transform 1 0 63020 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_685
timestamp 1644511149
transform 1 0 64124 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_697
timestamp 1644511149
transform 1 0 65228 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_709
timestamp 1644511149
transform 1 0 66332 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_721
timestamp 1644511149
transform 1 0 67436 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_727
timestamp 1644511149
transform 1 0 67988 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_729
timestamp 1644511149
transform 1 0 68172 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_7
timestamp 1644511149
transform 1 0 1748 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_19
timestamp 1644511149
transform 1 0 2852 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1644511149
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_29
timestamp 1644511149
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_41
timestamp 1644511149
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_53
timestamp 1644511149
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_65
timestamp 1644511149
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1644511149
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1644511149
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_85
timestamp 1644511149
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_97
timestamp 1644511149
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_109
timestamp 1644511149
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_121
timestamp 1644511149
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1644511149
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1644511149
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_100_141
timestamp 1644511149
transform 1 0 14076 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_146
timestamp 1644511149
transform 1 0 14536 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_150
timestamp 1644511149
transform 1 0 14904 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_156
timestamp 1644511149
transform 1 0 15456 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_168
timestamp 1644511149
transform 1 0 16560 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_175
timestamp 1644511149
transform 1 0 17204 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_183
timestamp 1644511149
transform 1 0 17940 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1644511149
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1644511149
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_197
timestamp 1644511149
transform 1 0 19228 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_205
timestamp 1644511149
transform 1 0 19964 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_212
timestamp 1644511149
transform 1 0 20608 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_220
timestamp 1644511149
transform 1 0 21344 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_229
timestamp 1644511149
transform 1 0 22172 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_241
timestamp 1644511149
transform 1 0 23276 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_249
timestamp 1644511149
transform 1 0 24012 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_253
timestamp 1644511149
transform 1 0 24380 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_261
timestamp 1644511149
transform 1 0 25116 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_269
timestamp 1644511149
transform 1 0 25852 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_288
timestamp 1644511149
transform 1 0 27600 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_296
timestamp 1644511149
transform 1 0 28336 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_309
timestamp 1644511149
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_321
timestamp 1644511149
transform 1 0 30636 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_100_339
timestamp 1644511149
transform 1 0 32292 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_347
timestamp 1644511149
transform 1 0 33028 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_353
timestamp 1644511149
transform 1 0 33580 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_360
timestamp 1644511149
transform 1 0 34224 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_365
timestamp 1644511149
transform 1 0 34684 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_373
timestamp 1644511149
transform 1 0 35420 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_381
timestamp 1644511149
transform 1 0 36156 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_398
timestamp 1644511149
transform 1 0 37720 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_406
timestamp 1644511149
transform 1 0 38456 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_414
timestamp 1644511149
transform 1 0 39192 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_100_421
timestamp 1644511149
transform 1 0 39836 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_429
timestamp 1644511149
transform 1 0 40572 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_100_447
timestamp 1644511149
transform 1 0 42228 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_455
timestamp 1644511149
transform 1 0 42964 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_472
timestamp 1644511149
transform 1 0 44528 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_477
timestamp 1644511149
transform 1 0 44988 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_483
timestamp 1644511149
transform 1 0 45540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_495
timestamp 1644511149
transform 1 0 46644 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_513
timestamp 1644511149
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1644511149
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1644511149
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_536
timestamp 1644511149
transform 1 0 50416 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_548
timestamp 1644511149
transform 1 0 51520 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_560
timestamp 1644511149
transform 1 0 52624 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_572
timestamp 1644511149
transform 1 0 53728 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_584
timestamp 1644511149
transform 1 0 54832 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_589
timestamp 1644511149
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_601
timestamp 1644511149
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_613
timestamp 1644511149
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_625
timestamp 1644511149
transform 1 0 58604 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_637
timestamp 1644511149
transform 1 0 59708 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_643
timestamp 1644511149
transform 1 0 60260 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_645
timestamp 1644511149
transform 1 0 60444 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_657
timestamp 1644511149
transform 1 0 61548 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_669
timestamp 1644511149
transform 1 0 62652 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_681
timestamp 1644511149
transform 1 0 63756 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_693
timestamp 1644511149
transform 1 0 64860 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_699
timestamp 1644511149
transform 1 0 65412 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_701
timestamp 1644511149
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_713
timestamp 1644511149
transform 1 0 66700 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_100_721
timestamp 1644511149
transform 1 0 67436 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_729
timestamp 1644511149
transform 1 0 68172 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_3
timestamp 1644511149
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_15
timestamp 1644511149
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_27
timestamp 1644511149
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_39
timestamp 1644511149
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_51
timestamp 1644511149
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1644511149
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1644511149
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1644511149
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_81
timestamp 1644511149
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_93
timestamp 1644511149
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_105
timestamp 1644511149
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1644511149
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_113
timestamp 1644511149
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_125
timestamp 1644511149
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_137
timestamp 1644511149
transform 1 0 13708 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_143
timestamp 1644511149
transform 1 0 14260 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_160
timestamp 1644511149
transform 1 0 15824 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_169
timestamp 1644511149
transform 1 0 16652 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_178
timestamp 1644511149
transform 1 0 17480 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_184
timestamp 1644511149
transform 1 0 18032 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_206
timestamp 1644511149
transform 1 0 20056 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_218
timestamp 1644511149
transform 1 0 21160 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_225
timestamp 1644511149
transform 1 0 21804 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_233
timestamp 1644511149
transform 1 0 22540 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_243
timestamp 1644511149
transform 1 0 23460 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_249
timestamp 1644511149
transform 1 0 24012 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_254
timestamp 1644511149
transform 1 0 24472 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_274
timestamp 1644511149
transform 1 0 26312 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_281
timestamp 1644511149
transform 1 0 26956 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_285
timestamp 1644511149
transform 1 0 27324 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_291
timestamp 1644511149
transform 1 0 27876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_303
timestamp 1644511149
transform 1 0 28980 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_311
timestamp 1644511149
transform 1 0 29716 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_318
timestamp 1644511149
transform 1 0 30360 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_326
timestamp 1644511149
transform 1 0 31096 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_334
timestamp 1644511149
transform 1 0 31832 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_345
timestamp 1644511149
transform 1 0 32844 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_353
timestamp 1644511149
transform 1 0 33580 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_375
timestamp 1644511149
transform 1 0 35604 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_384
timestamp 1644511149
transform 1 0 36432 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_101_398
timestamp 1644511149
transform 1 0 37720 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_406
timestamp 1644511149
transform 1 0 38456 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_413
timestamp 1644511149
transform 1 0 39100 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_421
timestamp 1644511149
transform 1 0 39836 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_433
timestamp 1644511149
transform 1 0 40940 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_438
timestamp 1644511149
transform 1 0 41400 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_446
timestamp 1644511149
transform 1 0 42136 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_449
timestamp 1644511149
transform 1 0 42412 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_456
timestamp 1644511149
transform 1 0 43056 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_468
timestamp 1644511149
transform 1 0 44160 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_480
timestamp 1644511149
transform 1 0 45264 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_492
timestamp 1644511149
transform 1 0 46368 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_505
timestamp 1644511149
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_517
timestamp 1644511149
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_529
timestamp 1644511149
transform 1 0 49772 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_541
timestamp 1644511149
transform 1 0 50876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_553
timestamp 1644511149
transform 1 0 51980 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1644511149
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_561
timestamp 1644511149
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_573
timestamp 1644511149
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_585
timestamp 1644511149
transform 1 0 54924 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_597
timestamp 1644511149
transform 1 0 56028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_609
timestamp 1644511149
transform 1 0 57132 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_615
timestamp 1644511149
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_617
timestamp 1644511149
transform 1 0 57868 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_629
timestamp 1644511149
transform 1 0 58972 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_641
timestamp 1644511149
transform 1 0 60076 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_653
timestamp 1644511149
transform 1 0 61180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_665
timestamp 1644511149
transform 1 0 62284 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_671
timestamp 1644511149
transform 1 0 62836 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_673
timestamp 1644511149
transform 1 0 63020 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_685
timestamp 1644511149
transform 1 0 64124 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_697
timestamp 1644511149
transform 1 0 65228 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_709
timestamp 1644511149
transform 1 0 66332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_724
timestamp 1644511149
transform 1 0 67712 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_729
timestamp 1644511149
transform 1 0 68172 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_3
timestamp 1644511149
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_15
timestamp 1644511149
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1644511149
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_29
timestamp 1644511149
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_41
timestamp 1644511149
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_53
timestamp 1644511149
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_65
timestamp 1644511149
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1644511149
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1644511149
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_85
timestamp 1644511149
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_97
timestamp 1644511149
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_109
timestamp 1644511149
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_121
timestamp 1644511149
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1644511149
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1644511149
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_141
timestamp 1644511149
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_153
timestamp 1644511149
transform 1 0 15180 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_102_163
timestamp 1644511149
transform 1 0 16100 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_183
timestamp 1644511149
transform 1 0 17940 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_195
timestamp 1644511149
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_102_197
timestamp 1644511149
transform 1 0 19228 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_102_208
timestamp 1644511149
transform 1 0 20240 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_102_218
timestamp 1644511149
transform 1 0 21160 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_102_230
timestamp 1644511149
transform 1 0 22264 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_102_248
timestamp 1644511149
transform 1 0 23920 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_274
timestamp 1644511149
transform 1 0 26312 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_294
timestamp 1644511149
transform 1 0 28152 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_102_306
timestamp 1644511149
transform 1 0 29256 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_102_309
timestamp 1644511149
transform 1 0 29532 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_313
timestamp 1644511149
transform 1 0 29900 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_102_333
timestamp 1644511149
transform 1 0 31740 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_339
timestamp 1644511149
transform 1 0 32292 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_356
timestamp 1644511149
transform 1 0 33856 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_102_381
timestamp 1644511149
transform 1 0 36156 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_102_390
timestamp 1644511149
transform 1 0 36984 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_402
timestamp 1644511149
transform 1 0 38088 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_406
timestamp 1644511149
transform 1 0 38456 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_410
timestamp 1644511149
transform 1 0 38824 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_102_418
timestamp 1644511149
transform 1 0 39560 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_102_421
timestamp 1644511149
transform 1 0 39836 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_433
timestamp 1644511149
transform 1 0 40940 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_445
timestamp 1644511149
transform 1 0 42044 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_457
timestamp 1644511149
transform 1 0 43148 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_102_465
timestamp 1644511149
transform 1 0 43884 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_102_470
timestamp 1644511149
transform 1 0 44344 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_102_493
timestamp 1644511149
transform 1 0 46460 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_505
timestamp 1644511149
transform 1 0 47564 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_517
timestamp 1644511149
transform 1 0 48668 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_102_529
timestamp 1644511149
transform 1 0 49772 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_102_533
timestamp 1644511149
transform 1 0 50140 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_545
timestamp 1644511149
transform 1 0 51244 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_557
timestamp 1644511149
transform 1 0 52348 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_569
timestamp 1644511149
transform 1 0 53452 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_581
timestamp 1644511149
transform 1 0 54556 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_587
timestamp 1644511149
transform 1 0 55108 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_589
timestamp 1644511149
transform 1 0 55292 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_601
timestamp 1644511149
transform 1 0 56396 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_613
timestamp 1644511149
transform 1 0 57500 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_625
timestamp 1644511149
transform 1 0 58604 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_637
timestamp 1644511149
transform 1 0 59708 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_643
timestamp 1644511149
transform 1 0 60260 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_645
timestamp 1644511149
transform 1 0 60444 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_657
timestamp 1644511149
transform 1 0 61548 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_669
timestamp 1644511149
transform 1 0 62652 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_681
timestamp 1644511149
transform 1 0 63756 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_693
timestamp 1644511149
transform 1 0 64860 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_699
timestamp 1644511149
transform 1 0 65412 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_102_701
timestamp 1644511149
transform 1 0 65596 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_707
timestamp 1644511149
transform 1 0 66148 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_729
timestamp 1644511149
transform 1 0 68172 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_3
timestamp 1644511149
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_15
timestamp 1644511149
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_27
timestamp 1644511149
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_39
timestamp 1644511149
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_51
timestamp 1644511149
transform 1 0 5796 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1644511149
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_57
timestamp 1644511149
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_69
timestamp 1644511149
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_81
timestamp 1644511149
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_93
timestamp 1644511149
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1644511149
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1644511149
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_113
timestamp 1644511149
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_125
timestamp 1644511149
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_137
timestamp 1644511149
transform 1 0 13708 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_103_143
timestamp 1644511149
transform 1 0 14260 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_147
timestamp 1644511149
transform 1 0 14628 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_153
timestamp 1644511149
transform 1 0 15180 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_103_165
timestamp 1644511149
transform 1 0 16284 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_103_169
timestamp 1644511149
transform 1 0 16652 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_175
timestamp 1644511149
transform 1 0 17204 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_187
timestamp 1644511149
transform 1 0 18308 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_103_211
timestamp 1644511149
transform 1 0 20516 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_220
timestamp 1644511149
transform 1 0 21344 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_103_241
timestamp 1644511149
transform 1 0 23276 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_103_249
timestamp 1644511149
transform 1 0 24012 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_103_255
timestamp 1644511149
transform 1 0 24564 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_261
timestamp 1644511149
transform 1 0 25116 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_267
timestamp 1644511149
transform 1 0 25668 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_271
timestamp 1644511149
transform 1 0 26036 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_276
timestamp 1644511149
transform 1 0 26496 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_103_281
timestamp 1644511149
transform 1 0 26956 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_103_286
timestamp 1644511149
transform 1 0 27416 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_290
timestamp 1644511149
transform 1 0 27784 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_312
timestamp 1644511149
transform 1 0 29808 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_103_320
timestamp 1644511149
transform 1 0 30544 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_103_329
timestamp 1644511149
transform 1 0 31372 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_335
timestamp 1644511149
transform 1 0 31924 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_103_343
timestamp 1644511149
transform 1 0 32660 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_103_351
timestamp 1644511149
transform 1 0 33396 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_103_356
timestamp 1644511149
transform 1 0 33856 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_368
timestamp 1644511149
transform 1 0 34960 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_380
timestamp 1644511149
transform 1 0 36064 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_396
timestamp 1644511149
transform 1 0 37536 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_400
timestamp 1644511149
transform 1 0 37904 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_405
timestamp 1644511149
transform 1 0 38364 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_409
timestamp 1644511149
transform 1 0 38732 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_416
timestamp 1644511149
transform 1 0 39376 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_424
timestamp 1644511149
transform 1 0 40112 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_432
timestamp 1644511149
transform 1 0 40848 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_103_442
timestamp 1644511149
transform 1 0 41768 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_103_449
timestamp 1644511149
transform 1 0 42412 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_103_457
timestamp 1644511149
transform 1 0 43148 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_465
timestamp 1644511149
transform 1 0 43884 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_474
timestamp 1644511149
transform 1 0 44712 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_486
timestamp 1644511149
transform 1 0 45816 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_498
timestamp 1644511149
transform 1 0 46920 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_103_505
timestamp 1644511149
transform 1 0 47564 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_517
timestamp 1644511149
transform 1 0 48668 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_529
timestamp 1644511149
transform 1 0 49772 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_541
timestamp 1644511149
transform 1 0 50876 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_553
timestamp 1644511149
transform 1 0 51980 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_559
timestamp 1644511149
transform 1 0 52532 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_561
timestamp 1644511149
transform 1 0 52716 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_573
timestamp 1644511149
transform 1 0 53820 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_585
timestamp 1644511149
transform 1 0 54924 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_597
timestamp 1644511149
transform 1 0 56028 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_609
timestamp 1644511149
transform 1 0 57132 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_615
timestamp 1644511149
transform 1 0 57684 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_617
timestamp 1644511149
transform 1 0 57868 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_629
timestamp 1644511149
transform 1 0 58972 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_641
timestamp 1644511149
transform 1 0 60076 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_653
timestamp 1644511149
transform 1 0 61180 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_665
timestamp 1644511149
transform 1 0 62284 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_671
timestamp 1644511149
transform 1 0 62836 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_673
timestamp 1644511149
transform 1 0 63020 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_685
timestamp 1644511149
transform 1 0 64124 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_697
timestamp 1644511149
transform 1 0 65228 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_709
timestamp 1644511149
transform 1 0 66332 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_724
timestamp 1644511149
transform 1 0 67712 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_729
timestamp 1644511149
transform 1 0 68172 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_104_3
timestamp 1644511149
transform 1 0 1380 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_104_12
timestamp 1644511149
transform 1 0 2208 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_104_24
timestamp 1644511149
transform 1 0 3312 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_104_29
timestamp 1644511149
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_41
timestamp 1644511149
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_53
timestamp 1644511149
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_65
timestamp 1644511149
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1644511149
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1644511149
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_85
timestamp 1644511149
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_97
timestamp 1644511149
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_109
timestamp 1644511149
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_121
timestamp 1644511149
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_133
timestamp 1644511149
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_139
timestamp 1644511149
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_157
timestamp 1644511149
transform 1 0 15548 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_169
timestamp 1644511149
transform 1 0 16652 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_180
timestamp 1644511149
transform 1 0 17664 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_104_192
timestamp 1644511149
transform 1 0 18768 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_201
timestamp 1644511149
transform 1 0 19596 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_104_208
timestamp 1644511149
transform 1 0 20240 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_220
timestamp 1644511149
transform 1 0 21344 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_224
timestamp 1644511149
transform 1 0 21712 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_236
timestamp 1644511149
transform 1 0 22816 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_104_248
timestamp 1644511149
transform 1 0 23920 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_104_253
timestamp 1644511149
transform 1 0 24380 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_261
timestamp 1644511149
transform 1 0 25116 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_265
timestamp 1644511149
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_277
timestamp 1644511149
transform 1 0 26588 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_289
timestamp 1644511149
transform 1 0 27692 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_301
timestamp 1644511149
transform 1 0 28796 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_307
timestamp 1644511149
transform 1 0 29348 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_314
timestamp 1644511149
transform 1 0 29992 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_104_326
timestamp 1644511149
transform 1 0 31096 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_104_336
timestamp 1644511149
transform 1 0 32016 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_348
timestamp 1644511149
transform 1 0 33120 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_104_360
timestamp 1644511149
transform 1 0 34224 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_104_365
timestamp 1644511149
transform 1 0 34684 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_104_383
timestamp 1644511149
transform 1 0 36340 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_391
timestamp 1644511149
transform 1 0 37076 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_397
timestamp 1644511149
transform 1 0 37628 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_104_405
timestamp 1644511149
transform 1 0 38364 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_104_415
timestamp 1644511149
transform 1 0 39284 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_104_419
timestamp 1644511149
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_428
timestamp 1644511149
transform 1 0 40480 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_104_448
timestamp 1644511149
transform 1 0 42320 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_454
timestamp 1644511149
transform 1 0 42872 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_459
timestamp 1644511149
transform 1 0 43332 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_104_471
timestamp 1644511149
transform 1 0 44436 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_104_475
timestamp 1644511149
transform 1 0 44804 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_477
timestamp 1644511149
transform 1 0 44988 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_489
timestamp 1644511149
transform 1 0 46092 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_501
timestamp 1644511149
transform 1 0 47196 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_513
timestamp 1644511149
transform 1 0 48300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_525
timestamp 1644511149
transform 1 0 49404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_531
timestamp 1644511149
transform 1 0 49956 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_533
timestamp 1644511149
transform 1 0 50140 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_545
timestamp 1644511149
transform 1 0 51244 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_557
timestamp 1644511149
transform 1 0 52348 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_569
timestamp 1644511149
transform 1 0 53452 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_581
timestamp 1644511149
transform 1 0 54556 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_587
timestamp 1644511149
transform 1 0 55108 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_589
timestamp 1644511149
transform 1 0 55292 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_601
timestamp 1644511149
transform 1 0 56396 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_613
timestamp 1644511149
transform 1 0 57500 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_625
timestamp 1644511149
transform 1 0 58604 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_637
timestamp 1644511149
transform 1 0 59708 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_643
timestamp 1644511149
transform 1 0 60260 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_645
timestamp 1644511149
transform 1 0 60444 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_657
timestamp 1644511149
transform 1 0 61548 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_669
timestamp 1644511149
transform 1 0 62652 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_681
timestamp 1644511149
transform 1 0 63756 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_693
timestamp 1644511149
transform 1 0 64860 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_699
timestamp 1644511149
transform 1 0 65412 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_701
timestamp 1644511149
transform 1 0 65596 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_713
timestamp 1644511149
transform 1 0 66700 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_725
timestamp 1644511149
transform 1 0 67804 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_105_3
timestamp 1644511149
transform 1 0 1380 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_105_27
timestamp 1644511149
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_39
timestamp 1644511149
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1644511149
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1644511149
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_57
timestamp 1644511149
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_69
timestamp 1644511149
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_81
timestamp 1644511149
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_93
timestamp 1644511149
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_105
timestamp 1644511149
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_111
timestamp 1644511149
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_113
timestamp 1644511149
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_125
timestamp 1644511149
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_137
timestamp 1644511149
transform 1 0 13708 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_105_148
timestamp 1644511149
transform 1 0 14720 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_156
timestamp 1644511149
transform 1 0 15456 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_105_162
timestamp 1644511149
transform 1 0 16008 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_105_174
timestamp 1644511149
transform 1 0 17112 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_105_182
timestamp 1644511149
transform 1 0 17848 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_211
timestamp 1644511149
transform 1 0 20516 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_223
timestamp 1644511149
transform 1 0 21620 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_225
timestamp 1644511149
transform 1 0 21804 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_232
timestamp 1644511149
transform 1 0 22448 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_105_252
timestamp 1644511149
transform 1 0 24288 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_105_260
timestamp 1644511149
transform 1 0 25024 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_266
timestamp 1644511149
transform 1 0 25576 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_105_278
timestamp 1644511149
transform 1 0 26680 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_105_297
timestamp 1644511149
transform 1 0 28428 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_305
timestamp 1644511149
transform 1 0 29164 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_105_323
timestamp 1644511149
transform 1 0 30820 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_335
timestamp 1644511149
transform 1 0 31924 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_105_337
timestamp 1644511149
transform 1 0 32108 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_346
timestamp 1644511149
transform 1 0 32936 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_105_354
timestamp 1644511149
transform 1 0 33672 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_376
timestamp 1644511149
transform 1 0 35696 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_105_386
timestamp 1644511149
transform 1 0 36616 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_105_409
timestamp 1644511149
transform 1 0 38732 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_415
timestamp 1644511149
transform 1 0 39284 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_426
timestamp 1644511149
transform 1 0 40296 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_442
timestamp 1644511149
transform 1 0 41768 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_105_449
timestamp 1644511149
transform 1 0 42412 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_105_462
timestamp 1644511149
transform 1 0 43608 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_469
timestamp 1644511149
transform 1 0 44252 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_481
timestamp 1644511149
transform 1 0 45356 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_493
timestamp 1644511149
transform 1 0 46460 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_105_501
timestamp 1644511149
transform 1 0 47196 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_105_505
timestamp 1644511149
transform 1 0 47564 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_517
timestamp 1644511149
transform 1 0 48668 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_529
timestamp 1644511149
transform 1 0 49772 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_541
timestamp 1644511149
transform 1 0 50876 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_553
timestamp 1644511149
transform 1 0 51980 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_559
timestamp 1644511149
transform 1 0 52532 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_561
timestamp 1644511149
transform 1 0 52716 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_573
timestamp 1644511149
transform 1 0 53820 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_585
timestamp 1644511149
transform 1 0 54924 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_597
timestamp 1644511149
transform 1 0 56028 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_609
timestamp 1644511149
transform 1 0 57132 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_615
timestamp 1644511149
transform 1 0 57684 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_617
timestamp 1644511149
transform 1 0 57868 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_629
timestamp 1644511149
transform 1 0 58972 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_641
timestamp 1644511149
transform 1 0 60076 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_653
timestamp 1644511149
transform 1 0 61180 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_665
timestamp 1644511149
transform 1 0 62284 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_671
timestamp 1644511149
transform 1 0 62836 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_673
timestamp 1644511149
transform 1 0 63020 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_685
timestamp 1644511149
transform 1 0 64124 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_697
timestamp 1644511149
transform 1 0 65228 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_709
timestamp 1644511149
transform 1 0 66332 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_105_717
timestamp 1644511149
transform 1 0 67068 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_724
timestamp 1644511149
transform 1 0 67712 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_729
timestamp 1644511149
transform 1 0 68172 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_3
timestamp 1644511149
transform 1 0 1380 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_9
timestamp 1644511149
transform 1 0 1932 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_21
timestamp 1644511149
transform 1 0 3036 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1644511149
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_29
timestamp 1644511149
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_41
timestamp 1644511149
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_53
timestamp 1644511149
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_65
timestamp 1644511149
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1644511149
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1644511149
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_85
timestamp 1644511149
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_97
timestamp 1644511149
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_109
timestamp 1644511149
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_121
timestamp 1644511149
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_133
timestamp 1644511149
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_139
timestamp 1644511149
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_141
timestamp 1644511149
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_153
timestamp 1644511149
transform 1 0 15180 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_173
timestamp 1644511149
transform 1 0 17020 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_182
timestamp 1644511149
transform 1 0 17848 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_106_194
timestamp 1644511149
transform 1 0 18952 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_106_197
timestamp 1644511149
transform 1 0 19228 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_209
timestamp 1644511149
transform 1 0 20332 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_213
timestamp 1644511149
transform 1 0 20700 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_235
timestamp 1644511149
transform 1 0 22724 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_243
timestamp 1644511149
transform 1 0 23460 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_248
timestamp 1644511149
transform 1 0 23920 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_269
timestamp 1644511149
transform 1 0 25852 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_277
timestamp 1644511149
transform 1 0 26588 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_106_304
timestamp 1644511149
transform 1 0 29072 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_312
timestamp 1644511149
transform 1 0 29808 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_106_324
timestamp 1644511149
transform 1 0 30912 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_106_334
timestamp 1644511149
transform 1 0 31832 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_342
timestamp 1644511149
transform 1 0 32568 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_359
timestamp 1644511149
transform 1 0 34132 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_363
timestamp 1644511149
transform 1 0 34500 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_106_365
timestamp 1644511149
transform 1 0 34684 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_371
timestamp 1644511149
transform 1 0 35236 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_375
timestamp 1644511149
transform 1 0 35604 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_387
timestamp 1644511149
transform 1 0 36708 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_399
timestamp 1644511149
transform 1 0 37812 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_407
timestamp 1644511149
transform 1 0 38548 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_106_415
timestamp 1644511149
transform 1 0 39284 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_419
timestamp 1644511149
transform 1 0 39652 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_425
timestamp 1644511149
transform 1 0 40204 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_437
timestamp 1644511149
transform 1 0 41308 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_449
timestamp 1644511149
transform 1 0 42412 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_453
timestamp 1644511149
transform 1 0 42780 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_106_470
timestamp 1644511149
transform 1 0 44344 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_106_477
timestamp 1644511149
transform 1 0 44988 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_489
timestamp 1644511149
transform 1 0 46092 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_501
timestamp 1644511149
transform 1 0 47196 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_513
timestamp 1644511149
transform 1 0 48300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_525
timestamp 1644511149
transform 1 0 49404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_531
timestamp 1644511149
transform 1 0 49956 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_533
timestamp 1644511149
transform 1 0 50140 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_545
timestamp 1644511149
transform 1 0 51244 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_557
timestamp 1644511149
transform 1 0 52348 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_569
timestamp 1644511149
transform 1 0 53452 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_581
timestamp 1644511149
transform 1 0 54556 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_587
timestamp 1644511149
transform 1 0 55108 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_589
timestamp 1644511149
transform 1 0 55292 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_601
timestamp 1644511149
transform 1 0 56396 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_613
timestamp 1644511149
transform 1 0 57500 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_625
timestamp 1644511149
transform 1 0 58604 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_637
timestamp 1644511149
transform 1 0 59708 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_643
timestamp 1644511149
transform 1 0 60260 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_645
timestamp 1644511149
transform 1 0 60444 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_657
timestamp 1644511149
transform 1 0 61548 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_669
timestamp 1644511149
transform 1 0 62652 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_681
timestamp 1644511149
transform 1 0 63756 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_693
timestamp 1644511149
transform 1 0 64860 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_699
timestamp 1644511149
transform 1 0 65412 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_701
timestamp 1644511149
transform 1 0 65596 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_713
timestamp 1644511149
transform 1 0 66700 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_106_722
timestamp 1644511149
transform 1 0 67528 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_729
timestamp 1644511149
transform 1 0 68172 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_3
timestamp 1644511149
transform 1 0 1380 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_13
timestamp 1644511149
transform 1 0 2300 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_25
timestamp 1644511149
transform 1 0 3404 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_37
timestamp 1644511149
transform 1 0 4508 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_49
timestamp 1644511149
transform 1 0 5612 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1644511149
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_57
timestamp 1644511149
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_69
timestamp 1644511149
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_81
timestamp 1644511149
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_93
timestamp 1644511149
transform 1 0 9660 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_105
timestamp 1644511149
transform 1 0 10764 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_111
timestamp 1644511149
transform 1 0 11316 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_113
timestamp 1644511149
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_125
timestamp 1644511149
transform 1 0 12604 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_137
timestamp 1644511149
transform 1 0 13708 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_149
timestamp 1644511149
transform 1 0 14812 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_164
timestamp 1644511149
transform 1 0 16192 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_107_169
timestamp 1644511149
transform 1 0 16652 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_107_193
timestamp 1644511149
transform 1 0 18860 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_199
timestamp 1644511149
transform 1 0 19412 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_203
timestamp 1644511149
transform 1 0 19780 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_215
timestamp 1644511149
transform 1 0 20884 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_223
timestamp 1644511149
transform 1 0 21620 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_225
timestamp 1644511149
transform 1 0 21804 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_107_234
timestamp 1644511149
transform 1 0 22632 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_242
timestamp 1644511149
transform 1 0 23368 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_246
timestamp 1644511149
transform 1 0 23736 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_107_258
timestamp 1644511149
transform 1 0 24840 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_107_262
timestamp 1644511149
transform 1 0 25208 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_270
timestamp 1644511149
transform 1 0 25944 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_276
timestamp 1644511149
transform 1 0 26496 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_107_281
timestamp 1644511149
transform 1 0 26956 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_289
timestamp 1644511149
transform 1 0 27692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_301
timestamp 1644511149
transform 1 0 28796 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_313
timestamp 1644511149
transform 1 0 29900 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_107_325
timestamp 1644511149
transform 1 0 31004 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_333
timestamp 1644511149
transform 1 0 31740 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_337
timestamp 1644511149
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_349
timestamp 1644511149
transform 1 0 33212 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_353
timestamp 1644511149
transform 1 0 33580 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_357
timestamp 1644511149
transform 1 0 33948 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_369
timestamp 1644511149
transform 1 0 35052 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_375
timestamp 1644511149
transform 1 0 35604 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_381
timestamp 1644511149
transform 1 0 36156 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_388
timestamp 1644511149
transform 1 0 36800 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_107_393
timestamp 1644511149
transform 1 0 37260 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_401
timestamp 1644511149
transform 1 0 37996 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_418
timestamp 1644511149
transform 1 0 39560 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_425
timestamp 1644511149
transform 1 0 40204 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_437
timestamp 1644511149
transform 1 0 41308 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_445
timestamp 1644511149
transform 1 0 42044 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_449
timestamp 1644511149
transform 1 0 42412 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_461
timestamp 1644511149
transform 1 0 43516 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_473
timestamp 1644511149
transform 1 0 44620 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_485
timestamp 1644511149
transform 1 0 45724 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_497
timestamp 1644511149
transform 1 0 46828 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_503
timestamp 1644511149
transform 1 0 47380 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_505
timestamp 1644511149
transform 1 0 47564 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_517
timestamp 1644511149
transform 1 0 48668 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_529
timestamp 1644511149
transform 1 0 49772 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_541
timestamp 1644511149
transform 1 0 50876 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_553
timestamp 1644511149
transform 1 0 51980 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_559
timestamp 1644511149
transform 1 0 52532 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_561
timestamp 1644511149
transform 1 0 52716 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_573
timestamp 1644511149
transform 1 0 53820 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_585
timestamp 1644511149
transform 1 0 54924 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_597
timestamp 1644511149
transform 1 0 56028 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_609
timestamp 1644511149
transform 1 0 57132 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_615
timestamp 1644511149
transform 1 0 57684 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_617
timestamp 1644511149
transform 1 0 57868 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_629
timestamp 1644511149
transform 1 0 58972 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_641
timestamp 1644511149
transform 1 0 60076 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_653
timestamp 1644511149
transform 1 0 61180 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_665
timestamp 1644511149
transform 1 0 62284 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_671
timestamp 1644511149
transform 1 0 62836 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_673
timestamp 1644511149
transform 1 0 63020 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_685
timestamp 1644511149
transform 1 0 64124 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_697
timestamp 1644511149
transform 1 0 65228 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_107_724
timestamp 1644511149
transform 1 0 67712 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_729
timestamp 1644511149
transform 1 0 68172 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_108_3
timestamp 1644511149
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_15
timestamp 1644511149
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1644511149
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_29
timestamp 1644511149
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_41
timestamp 1644511149
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_53
timestamp 1644511149
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_65
timestamp 1644511149
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1644511149
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1644511149
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_85
timestamp 1644511149
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_97
timestamp 1644511149
transform 1 0 10028 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_109
timestamp 1644511149
transform 1 0 11132 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_121
timestamp 1644511149
transform 1 0 12236 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_133
timestamp 1644511149
transform 1 0 13340 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_139
timestamp 1644511149
transform 1 0 13892 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_141
timestamp 1644511149
transform 1 0 14076 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_153
timestamp 1644511149
transform 1 0 15180 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_165
timestamp 1644511149
transform 1 0 16284 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_177
timestamp 1644511149
transform 1 0 17388 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_189
timestamp 1644511149
transform 1 0 18492 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_195
timestamp 1644511149
transform 1 0 19044 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_197
timestamp 1644511149
transform 1 0 19228 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_204
timestamp 1644511149
transform 1 0 19872 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_208
timestamp 1644511149
transform 1 0 20240 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_214
timestamp 1644511149
transform 1 0 20792 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_234
timestamp 1644511149
transform 1 0 22632 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_242
timestamp 1644511149
transform 1 0 23368 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_246
timestamp 1644511149
transform 1 0 23736 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_108_265
timestamp 1644511149
transform 1 0 25484 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_273
timestamp 1644511149
transform 1 0 26220 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_108_278
timestamp 1644511149
transform 1 0 26680 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_284
timestamp 1644511149
transform 1 0 27232 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_290
timestamp 1644511149
transform 1 0 27784 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_294
timestamp 1644511149
transform 1 0 28152 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_300
timestamp 1644511149
transform 1 0 28704 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_108_309
timestamp 1644511149
transform 1 0 29532 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_108_317
timestamp 1644511149
transform 1 0 30268 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_328
timestamp 1644511149
transform 1 0 31280 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_108_348
timestamp 1644511149
transform 1 0 33120 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_108_360
timestamp 1644511149
transform 1 0 34224 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_365
timestamp 1644511149
transform 1 0 34684 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_370
timestamp 1644511149
transform 1 0 35144 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_108_384
timestamp 1644511149
transform 1 0 36432 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_404
timestamp 1644511149
transform 1 0 38272 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_412
timestamp 1644511149
transform 1 0 39008 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_437
timestamp 1644511149
transform 1 0 41308 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_449
timestamp 1644511149
transform 1 0 42412 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_461
timestamp 1644511149
transform 1 0 43516 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_108_473
timestamp 1644511149
transform 1 0 44620 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_477
timestamp 1644511149
transform 1 0 44988 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_489
timestamp 1644511149
transform 1 0 46092 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_501
timestamp 1644511149
transform 1 0 47196 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_513
timestamp 1644511149
transform 1 0 48300 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_525
timestamp 1644511149
transform 1 0 49404 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_531
timestamp 1644511149
transform 1 0 49956 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_533
timestamp 1644511149
transform 1 0 50140 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_545
timestamp 1644511149
transform 1 0 51244 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_557
timestamp 1644511149
transform 1 0 52348 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_569
timestamp 1644511149
transform 1 0 53452 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_581
timestamp 1644511149
transform 1 0 54556 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_587
timestamp 1644511149
transform 1 0 55108 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_589
timestamp 1644511149
transform 1 0 55292 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_601
timestamp 1644511149
transform 1 0 56396 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_613
timestamp 1644511149
transform 1 0 57500 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_625
timestamp 1644511149
transform 1 0 58604 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_637
timestamp 1644511149
transform 1 0 59708 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_643
timestamp 1644511149
transform 1 0 60260 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_645
timestamp 1644511149
transform 1 0 60444 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_657
timestamp 1644511149
transform 1 0 61548 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_669
timestamp 1644511149
transform 1 0 62652 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_681
timestamp 1644511149
transform 1 0 63756 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_693
timestamp 1644511149
transform 1 0 64860 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_699
timestamp 1644511149
transform 1 0 65412 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_701
timestamp 1644511149
transform 1 0 65596 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_713
timestamp 1644511149
transform 1 0 66700 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_721
timestamp 1644511149
transform 1 0 67436 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_725
timestamp 1644511149
transform 1 0 67804 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_3
timestamp 1644511149
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_15
timestamp 1644511149
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_27
timestamp 1644511149
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_39
timestamp 1644511149
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_51
timestamp 1644511149
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1644511149
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_57
timestamp 1644511149
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_69
timestamp 1644511149
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_81
timestamp 1644511149
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_93
timestamp 1644511149
transform 1 0 9660 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_105
timestamp 1644511149
transform 1 0 10764 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_111
timestamp 1644511149
transform 1 0 11316 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_113
timestamp 1644511149
transform 1 0 11500 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_125
timestamp 1644511149
transform 1 0 12604 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_137
timestamp 1644511149
transform 1 0 13708 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_149
timestamp 1644511149
transform 1 0 14812 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_161
timestamp 1644511149
transform 1 0 15916 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_167
timestamp 1644511149
transform 1 0 16468 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_169
timestamp 1644511149
transform 1 0 16652 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_181
timestamp 1644511149
transform 1 0 17756 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_193
timestamp 1644511149
transform 1 0 18860 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_213
timestamp 1644511149
transform 1 0 20700 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_220
timestamp 1644511149
transform 1 0 21344 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_109_229
timestamp 1644511149
transform 1 0 22172 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_109_256
timestamp 1644511149
transform 1 0 24656 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_266
timestamp 1644511149
transform 1 0 25576 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_109_274
timestamp 1644511149
transform 1 0 26312 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_109_281
timestamp 1644511149
transform 1 0 26956 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_109_303
timestamp 1644511149
transform 1 0 28980 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_309
timestamp 1644511149
transform 1 0 29532 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_109_326
timestamp 1644511149
transform 1 0 31096 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_334
timestamp 1644511149
transform 1 0 31832 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_109_337
timestamp 1644511149
transform 1 0 32108 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_349
timestamp 1644511149
transform 1 0 33212 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_109_367
timestamp 1644511149
transform 1 0 34868 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_375
timestamp 1644511149
transform 1 0 35604 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_109_384
timestamp 1644511149
transform 1 0 36432 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_393
timestamp 1644511149
transform 1 0 37260 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_405
timestamp 1644511149
transform 1 0 38364 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_417
timestamp 1644511149
transform 1 0 39468 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_429
timestamp 1644511149
transform 1 0 40572 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_441
timestamp 1644511149
transform 1 0 41676 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_447
timestamp 1644511149
transform 1 0 42228 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_449
timestamp 1644511149
transform 1 0 42412 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_461
timestamp 1644511149
transform 1 0 43516 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_473
timestamp 1644511149
transform 1 0 44620 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_485
timestamp 1644511149
transform 1 0 45724 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_497
timestamp 1644511149
transform 1 0 46828 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_503
timestamp 1644511149
transform 1 0 47380 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_505
timestamp 1644511149
transform 1 0 47564 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_517
timestamp 1644511149
transform 1 0 48668 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_529
timestamp 1644511149
transform 1 0 49772 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_541
timestamp 1644511149
transform 1 0 50876 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_553
timestamp 1644511149
transform 1 0 51980 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_559
timestamp 1644511149
transform 1 0 52532 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_561
timestamp 1644511149
transform 1 0 52716 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_573
timestamp 1644511149
transform 1 0 53820 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_585
timestamp 1644511149
transform 1 0 54924 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_597
timestamp 1644511149
transform 1 0 56028 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_609
timestamp 1644511149
transform 1 0 57132 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_615
timestamp 1644511149
transform 1 0 57684 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_617
timestamp 1644511149
transform 1 0 57868 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_629
timestamp 1644511149
transform 1 0 58972 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_641
timestamp 1644511149
transform 1 0 60076 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_653
timestamp 1644511149
transform 1 0 61180 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_665
timestamp 1644511149
transform 1 0 62284 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_671
timestamp 1644511149
transform 1 0 62836 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_673
timestamp 1644511149
transform 1 0 63020 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_685
timestamp 1644511149
transform 1 0 64124 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_697
timestamp 1644511149
transform 1 0 65228 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_109_724
timestamp 1644511149
transform 1 0 67712 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_729
timestamp 1644511149
transform 1 0 68172 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_110_3
timestamp 1644511149
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_15
timestamp 1644511149
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1644511149
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_29
timestamp 1644511149
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_41
timestamp 1644511149
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_53
timestamp 1644511149
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_65
timestamp 1644511149
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1644511149
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1644511149
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_85
timestamp 1644511149
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_97
timestamp 1644511149
transform 1 0 10028 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_109
timestamp 1644511149
transform 1 0 11132 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_121
timestamp 1644511149
transform 1 0 12236 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_133
timestamp 1644511149
transform 1 0 13340 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_139
timestamp 1644511149
transform 1 0 13892 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_141
timestamp 1644511149
transform 1 0 14076 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_153
timestamp 1644511149
transform 1 0 15180 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_165
timestamp 1644511149
transform 1 0 16284 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_177
timestamp 1644511149
transform 1 0 17388 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_189
timestamp 1644511149
transform 1 0 18492 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_195
timestamp 1644511149
transform 1 0 19044 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_110_197
timestamp 1644511149
transform 1 0 19228 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_201
timestamp 1644511149
transform 1 0 19596 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_206
timestamp 1644511149
transform 1 0 20056 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_218
timestamp 1644511149
transform 1 0 21160 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_110_230
timestamp 1644511149
transform 1 0 22264 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_110_248
timestamp 1644511149
transform 1 0 23920 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_269
timestamp 1644511149
transform 1 0 25852 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_289
timestamp 1644511149
transform 1 0 27692 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_297
timestamp 1644511149
transform 1 0 28428 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_304
timestamp 1644511149
transform 1 0 29072 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_110_309
timestamp 1644511149
transform 1 0 29532 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_110_314
timestamp 1644511149
transform 1 0 29992 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_110_339
timestamp 1644511149
transform 1 0 32292 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_350
timestamp 1644511149
transform 1 0 33304 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_110_362
timestamp 1644511149
transform 1 0 34408 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_110_365
timestamp 1644511149
transform 1 0 34684 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_110_375
timestamp 1644511149
transform 1 0 35604 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_387
timestamp 1644511149
transform 1 0 36708 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_110_395
timestamp 1644511149
transform 1 0 37444 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_406
timestamp 1644511149
transform 1 0 38456 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_110_418
timestamp 1644511149
transform 1 0 39560 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_110_421
timestamp 1644511149
transform 1 0 39836 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_433
timestamp 1644511149
transform 1 0 40940 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_445
timestamp 1644511149
transform 1 0 42044 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_457
timestamp 1644511149
transform 1 0 43148 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_469
timestamp 1644511149
transform 1 0 44252 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_475
timestamp 1644511149
transform 1 0 44804 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_477
timestamp 1644511149
transform 1 0 44988 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_489
timestamp 1644511149
transform 1 0 46092 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_501
timestamp 1644511149
transform 1 0 47196 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_513
timestamp 1644511149
transform 1 0 48300 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_525
timestamp 1644511149
transform 1 0 49404 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_531
timestamp 1644511149
transform 1 0 49956 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_533
timestamp 1644511149
transform 1 0 50140 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_545
timestamp 1644511149
transform 1 0 51244 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_557
timestamp 1644511149
transform 1 0 52348 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_569
timestamp 1644511149
transform 1 0 53452 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_581
timestamp 1644511149
transform 1 0 54556 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_587
timestamp 1644511149
transform 1 0 55108 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_589
timestamp 1644511149
transform 1 0 55292 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_601
timestamp 1644511149
transform 1 0 56396 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_613
timestamp 1644511149
transform 1 0 57500 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_625
timestamp 1644511149
transform 1 0 58604 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_637
timestamp 1644511149
transform 1 0 59708 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_643
timestamp 1644511149
transform 1 0 60260 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_645
timestamp 1644511149
transform 1 0 60444 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_657
timestamp 1644511149
transform 1 0 61548 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_669
timestamp 1644511149
transform 1 0 62652 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_681
timestamp 1644511149
transform 1 0 63756 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_693
timestamp 1644511149
transform 1 0 64860 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_699
timestamp 1644511149
transform 1 0 65412 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_701
timestamp 1644511149
transform 1 0 65596 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_713
timestamp 1644511149
transform 1 0 66700 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_110_721
timestamp 1644511149
transform 1 0 67436 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_110_727
timestamp 1644511149
transform 1 0 67988 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_111_3
timestamp 1644511149
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_15
timestamp 1644511149
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_27
timestamp 1644511149
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_39
timestamp 1644511149
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_51
timestamp 1644511149
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1644511149
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_57
timestamp 1644511149
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_69
timestamp 1644511149
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_81
timestamp 1644511149
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_93
timestamp 1644511149
transform 1 0 9660 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_105
timestamp 1644511149
transform 1 0 10764 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_111
timestamp 1644511149
transform 1 0 11316 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_113
timestamp 1644511149
transform 1 0 11500 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_125
timestamp 1644511149
transform 1 0 12604 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_137
timestamp 1644511149
transform 1 0 13708 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_149
timestamp 1644511149
transform 1 0 14812 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_161
timestamp 1644511149
transform 1 0 15916 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_167
timestamp 1644511149
transform 1 0 16468 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_169
timestamp 1644511149
transform 1 0 16652 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_181
timestamp 1644511149
transform 1 0 17756 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_193
timestamp 1644511149
transform 1 0 18860 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_205
timestamp 1644511149
transform 1 0 19964 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_217
timestamp 1644511149
transform 1 0 21068 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_223
timestamp 1644511149
transform 1 0 21620 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_225
timestamp 1644511149
transform 1 0 21804 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_111_237
timestamp 1644511149
transform 1 0 22908 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_111_244
timestamp 1644511149
transform 1 0 23552 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_111_264
timestamp 1644511149
transform 1 0 25392 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_276
timestamp 1644511149
transform 1 0 26496 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_111_281
timestamp 1644511149
transform 1 0 26956 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_293
timestamp 1644511149
transform 1 0 28060 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_111_300
timestamp 1644511149
transform 1 0 28704 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_111_325
timestamp 1644511149
transform 1 0 31004 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_111_333
timestamp 1644511149
transform 1 0 31740 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_111_337
timestamp 1644511149
transform 1 0 32108 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_111_345
timestamp 1644511149
transform 1 0 32844 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_111_367
timestamp 1644511149
transform 1 0 34868 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_371
timestamp 1644511149
transform 1 0 35236 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_111_377
timestamp 1644511149
transform 1 0 35788 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_111_387
timestamp 1644511149
transform 1 0 36708 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_391
timestamp 1644511149
transform 1 0 37076 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_111_393
timestamp 1644511149
transform 1 0 37260 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_111_400
timestamp 1644511149
transform 1 0 37904 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_111_420
timestamp 1644511149
transform 1 0 39744 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_432
timestamp 1644511149
transform 1 0 40848 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_444
timestamp 1644511149
transform 1 0 41952 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_111_449
timestamp 1644511149
transform 1 0 42412 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_461
timestamp 1644511149
transform 1 0 43516 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_473
timestamp 1644511149
transform 1 0 44620 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_485
timestamp 1644511149
transform 1 0 45724 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_497
timestamp 1644511149
transform 1 0 46828 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_503
timestamp 1644511149
transform 1 0 47380 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_505
timestamp 1644511149
transform 1 0 47564 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_517
timestamp 1644511149
transform 1 0 48668 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_529
timestamp 1644511149
transform 1 0 49772 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_541
timestamp 1644511149
transform 1 0 50876 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_553
timestamp 1644511149
transform 1 0 51980 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_559
timestamp 1644511149
transform 1 0 52532 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_561
timestamp 1644511149
transform 1 0 52716 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_573
timestamp 1644511149
transform 1 0 53820 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_585
timestamp 1644511149
transform 1 0 54924 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_597
timestamp 1644511149
transform 1 0 56028 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_609
timestamp 1644511149
transform 1 0 57132 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_615
timestamp 1644511149
transform 1 0 57684 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_617
timestamp 1644511149
transform 1 0 57868 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_629
timestamp 1644511149
transform 1 0 58972 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_641
timestamp 1644511149
transform 1 0 60076 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_653
timestamp 1644511149
transform 1 0 61180 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_665
timestamp 1644511149
transform 1 0 62284 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_671
timestamp 1644511149
transform 1 0 62836 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_673
timestamp 1644511149
transform 1 0 63020 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_685
timestamp 1644511149
transform 1 0 64124 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_697
timestamp 1644511149
transform 1 0 65228 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_709
timestamp 1644511149
transform 1 0 66332 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_724
timestamp 1644511149
transform 1 0 67712 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_111_729
timestamp 1644511149
transform 1 0 68172 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_112_9
timestamp 1644511149
transform 1 0 1932 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_21
timestamp 1644511149
transform 1 0 3036 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1644511149
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_29
timestamp 1644511149
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_41
timestamp 1644511149
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_53
timestamp 1644511149
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_65
timestamp 1644511149
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_77
timestamp 1644511149
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_83
timestamp 1644511149
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_85
timestamp 1644511149
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_97
timestamp 1644511149
transform 1 0 10028 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_109
timestamp 1644511149
transform 1 0 11132 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_121
timestamp 1644511149
transform 1 0 12236 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_133
timestamp 1644511149
transform 1 0 13340 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_139
timestamp 1644511149
transform 1 0 13892 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_141
timestamp 1644511149
transform 1 0 14076 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_153
timestamp 1644511149
transform 1 0 15180 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_165
timestamp 1644511149
transform 1 0 16284 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_177
timestamp 1644511149
transform 1 0 17388 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_189
timestamp 1644511149
transform 1 0 18492 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_195
timestamp 1644511149
transform 1 0 19044 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_197
timestamp 1644511149
transform 1 0 19228 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_209
timestamp 1644511149
transform 1 0 20332 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_221
timestamp 1644511149
transform 1 0 21436 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_233
timestamp 1644511149
transform 1 0 22540 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_245
timestamp 1644511149
transform 1 0 23644 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_251
timestamp 1644511149
transform 1 0 24196 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_262
timestamp 1644511149
transform 1 0 25208 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_274
timestamp 1644511149
transform 1 0 26312 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_286
timestamp 1644511149
transform 1 0 27416 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_298
timestamp 1644511149
transform 1 0 28520 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_112_306
timestamp 1644511149
transform 1 0 29256 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_112_309
timestamp 1644511149
transform 1 0 29532 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_321
timestamp 1644511149
transform 1 0 30636 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_333
timestamp 1644511149
transform 1 0 31740 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_345
timestamp 1644511149
transform 1 0 32844 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_357
timestamp 1644511149
transform 1 0 33948 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_363
timestamp 1644511149
transform 1 0 34500 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_112_368
timestamp 1644511149
transform 1 0 34960 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_374
timestamp 1644511149
transform 1 0 35512 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_112_382
timestamp 1644511149
transform 1 0 36248 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_112_386
timestamp 1644511149
transform 1 0 36616 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_394
timestamp 1644511149
transform 1 0 37352 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_406
timestamp 1644511149
transform 1 0 38456 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_112_418
timestamp 1644511149
transform 1 0 39560 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_112_421
timestamp 1644511149
transform 1 0 39836 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_433
timestamp 1644511149
transform 1 0 40940 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_445
timestamp 1644511149
transform 1 0 42044 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_457
timestamp 1644511149
transform 1 0 43148 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_469
timestamp 1644511149
transform 1 0 44252 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_475
timestamp 1644511149
transform 1 0 44804 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_477
timestamp 1644511149
transform 1 0 44988 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_489
timestamp 1644511149
transform 1 0 46092 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_501
timestamp 1644511149
transform 1 0 47196 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_513
timestamp 1644511149
transform 1 0 48300 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_525
timestamp 1644511149
transform 1 0 49404 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_531
timestamp 1644511149
transform 1 0 49956 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_533
timestamp 1644511149
transform 1 0 50140 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_545
timestamp 1644511149
transform 1 0 51244 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_557
timestamp 1644511149
transform 1 0 52348 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_569
timestamp 1644511149
transform 1 0 53452 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_581
timestamp 1644511149
transform 1 0 54556 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_587
timestamp 1644511149
transform 1 0 55108 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_589
timestamp 1644511149
transform 1 0 55292 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_601
timestamp 1644511149
transform 1 0 56396 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_613
timestamp 1644511149
transform 1 0 57500 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_625
timestamp 1644511149
transform 1 0 58604 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_637
timestamp 1644511149
transform 1 0 59708 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_643
timestamp 1644511149
transform 1 0 60260 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_645
timestamp 1644511149
transform 1 0 60444 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_657
timestamp 1644511149
transform 1 0 61548 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_669
timestamp 1644511149
transform 1 0 62652 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_681
timestamp 1644511149
transform 1 0 63756 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_693
timestamp 1644511149
transform 1 0 64860 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_699
timestamp 1644511149
transform 1 0 65412 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_112_701
timestamp 1644511149
transform 1 0 65596 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_707
timestamp 1644511149
transform 1 0 66148 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_112_729
timestamp 1644511149
transform 1 0 68172 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_113_3
timestamp 1644511149
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_15
timestamp 1644511149
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_27
timestamp 1644511149
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_39
timestamp 1644511149
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1644511149
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1644511149
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_57
timestamp 1644511149
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_69
timestamp 1644511149
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_81
timestamp 1644511149
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_93
timestamp 1644511149
transform 1 0 9660 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_105
timestamp 1644511149
transform 1 0 10764 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_111
timestamp 1644511149
transform 1 0 11316 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_113
timestamp 1644511149
transform 1 0 11500 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_125
timestamp 1644511149
transform 1 0 12604 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_137
timestamp 1644511149
transform 1 0 13708 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_149
timestamp 1644511149
transform 1 0 14812 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_161
timestamp 1644511149
transform 1 0 15916 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_167
timestamp 1644511149
transform 1 0 16468 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_169
timestamp 1644511149
transform 1 0 16652 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_181
timestamp 1644511149
transform 1 0 17756 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_193
timestamp 1644511149
transform 1 0 18860 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_205
timestamp 1644511149
transform 1 0 19964 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_217
timestamp 1644511149
transform 1 0 21068 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_223
timestamp 1644511149
transform 1 0 21620 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_225
timestamp 1644511149
transform 1 0 21804 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_237
timestamp 1644511149
transform 1 0 22908 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_249
timestamp 1644511149
transform 1 0 24012 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_261
timestamp 1644511149
transform 1 0 25116 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_273
timestamp 1644511149
transform 1 0 26220 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_279
timestamp 1644511149
transform 1 0 26772 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_281
timestamp 1644511149
transform 1 0 26956 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_293
timestamp 1644511149
transform 1 0 28060 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_305
timestamp 1644511149
transform 1 0 29164 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_317
timestamp 1644511149
transform 1 0 30268 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_329
timestamp 1644511149
transform 1 0 31372 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_335
timestamp 1644511149
transform 1 0 31924 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_337
timestamp 1644511149
transform 1 0 32108 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_349
timestamp 1644511149
transform 1 0 33212 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_113_373
timestamp 1644511149
transform 1 0 35420 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_113_381
timestamp 1644511149
transform 1 0 36156 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_113_388
timestamp 1644511149
transform 1 0 36800 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_113_393
timestamp 1644511149
transform 1 0 37260 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_113_402
timestamp 1644511149
transform 1 0 38088 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_414
timestamp 1644511149
transform 1 0 39192 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_426
timestamp 1644511149
transform 1 0 40296 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_438
timestamp 1644511149
transform 1 0 41400 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_113_446
timestamp 1644511149
transform 1 0 42136 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_113_449
timestamp 1644511149
transform 1 0 42412 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_461
timestamp 1644511149
transform 1 0 43516 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_473
timestamp 1644511149
transform 1 0 44620 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_485
timestamp 1644511149
transform 1 0 45724 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_497
timestamp 1644511149
transform 1 0 46828 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_503
timestamp 1644511149
transform 1 0 47380 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_505
timestamp 1644511149
transform 1 0 47564 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_517
timestamp 1644511149
transform 1 0 48668 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_529
timestamp 1644511149
transform 1 0 49772 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_541
timestamp 1644511149
transform 1 0 50876 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_553
timestamp 1644511149
transform 1 0 51980 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_559
timestamp 1644511149
transform 1 0 52532 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_561
timestamp 1644511149
transform 1 0 52716 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_573
timestamp 1644511149
transform 1 0 53820 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_585
timestamp 1644511149
transform 1 0 54924 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_597
timestamp 1644511149
transform 1 0 56028 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_609
timestamp 1644511149
transform 1 0 57132 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_615
timestamp 1644511149
transform 1 0 57684 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_617
timestamp 1644511149
transform 1 0 57868 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_629
timestamp 1644511149
transform 1 0 58972 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_641
timestamp 1644511149
transform 1 0 60076 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_653
timestamp 1644511149
transform 1 0 61180 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_665
timestamp 1644511149
transform 1 0 62284 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_671
timestamp 1644511149
transform 1 0 62836 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_673
timestamp 1644511149
transform 1 0 63020 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_685
timestamp 1644511149
transform 1 0 64124 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_697
timestamp 1644511149
transform 1 0 65228 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_709
timestamp 1644511149
transform 1 0 66332 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_724
timestamp 1644511149
transform 1 0 67712 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_729
timestamp 1644511149
transform 1 0 68172 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_3
timestamp 1644511149
transform 1 0 1380 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_114_10
timestamp 1644511149
transform 1 0 2024 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_22
timestamp 1644511149
transform 1 0 3128 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_114_29
timestamp 1644511149
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_41
timestamp 1644511149
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_53
timestamp 1644511149
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_65
timestamp 1644511149
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1644511149
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1644511149
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_85
timestamp 1644511149
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_97
timestamp 1644511149
transform 1 0 10028 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_109
timestamp 1644511149
transform 1 0 11132 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_121
timestamp 1644511149
transform 1 0 12236 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_133
timestamp 1644511149
transform 1 0 13340 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_139
timestamp 1644511149
transform 1 0 13892 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_141
timestamp 1644511149
transform 1 0 14076 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_153
timestamp 1644511149
transform 1 0 15180 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_165
timestamp 1644511149
transform 1 0 16284 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_177
timestamp 1644511149
transform 1 0 17388 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_189
timestamp 1644511149
transform 1 0 18492 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_195
timestamp 1644511149
transform 1 0 19044 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_197
timestamp 1644511149
transform 1 0 19228 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_209
timestamp 1644511149
transform 1 0 20332 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_221
timestamp 1644511149
transform 1 0 21436 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_233
timestamp 1644511149
transform 1 0 22540 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_245
timestamp 1644511149
transform 1 0 23644 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_251
timestamp 1644511149
transform 1 0 24196 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_253
timestamp 1644511149
transform 1 0 24380 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_265
timestamp 1644511149
transform 1 0 25484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_277
timestamp 1644511149
transform 1 0 26588 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_289
timestamp 1644511149
transform 1 0 27692 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_301
timestamp 1644511149
transform 1 0 28796 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_307
timestamp 1644511149
transform 1 0 29348 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_309
timestamp 1644511149
transform 1 0 29532 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_321
timestamp 1644511149
transform 1 0 30636 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_333
timestamp 1644511149
transform 1 0 31740 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_345
timestamp 1644511149
transform 1 0 32844 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_357
timestamp 1644511149
transform 1 0 33948 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_363
timestamp 1644511149
transform 1 0 34500 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_365
timestamp 1644511149
transform 1 0 34684 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_114_377
timestamp 1644511149
transform 1 0 35788 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_385
timestamp 1644511149
transform 1 0 36524 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_396
timestamp 1644511149
transform 1 0 37536 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_416
timestamp 1644511149
transform 1 0 39376 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_114_421
timestamp 1644511149
transform 1 0 39836 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_433
timestamp 1644511149
transform 1 0 40940 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_445
timestamp 1644511149
transform 1 0 42044 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_457
timestamp 1644511149
transform 1 0 43148 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_469
timestamp 1644511149
transform 1 0 44252 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_475
timestamp 1644511149
transform 1 0 44804 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_477
timestamp 1644511149
transform 1 0 44988 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_489
timestamp 1644511149
transform 1 0 46092 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_501
timestamp 1644511149
transform 1 0 47196 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_513
timestamp 1644511149
transform 1 0 48300 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_525
timestamp 1644511149
transform 1 0 49404 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_531
timestamp 1644511149
transform 1 0 49956 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_533
timestamp 1644511149
transform 1 0 50140 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_545
timestamp 1644511149
transform 1 0 51244 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_557
timestamp 1644511149
transform 1 0 52348 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_569
timestamp 1644511149
transform 1 0 53452 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_581
timestamp 1644511149
transform 1 0 54556 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_587
timestamp 1644511149
transform 1 0 55108 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_589
timestamp 1644511149
transform 1 0 55292 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_601
timestamp 1644511149
transform 1 0 56396 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_613
timestamp 1644511149
transform 1 0 57500 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_625
timestamp 1644511149
transform 1 0 58604 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_637
timestamp 1644511149
transform 1 0 59708 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_643
timestamp 1644511149
transform 1 0 60260 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_645
timestamp 1644511149
transform 1 0 60444 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_657
timestamp 1644511149
transform 1 0 61548 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_669
timestamp 1644511149
transform 1 0 62652 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_681
timestamp 1644511149
transform 1 0 63756 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_693
timestamp 1644511149
transform 1 0 64860 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_699
timestamp 1644511149
transform 1 0 65412 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_701
timestamp 1644511149
transform 1 0 65596 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_713
timestamp 1644511149
transform 1 0 66700 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_725
timestamp 1644511149
transform 1 0 67804 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_115_3
timestamp 1644511149
transform 1 0 1380 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_28
timestamp 1644511149
transform 1 0 3680 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_115_38
timestamp 1644511149
transform 1 0 4600 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_50
timestamp 1644511149
transform 1 0 5704 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_115_57
timestamp 1644511149
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_69
timestamp 1644511149
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_81
timestamp 1644511149
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_93
timestamp 1644511149
transform 1 0 9660 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_105
timestamp 1644511149
transform 1 0 10764 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_111
timestamp 1644511149
transform 1 0 11316 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_113
timestamp 1644511149
transform 1 0 11500 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_125
timestamp 1644511149
transform 1 0 12604 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_137
timestamp 1644511149
transform 1 0 13708 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_149
timestamp 1644511149
transform 1 0 14812 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_161
timestamp 1644511149
transform 1 0 15916 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_167
timestamp 1644511149
transform 1 0 16468 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_169
timestamp 1644511149
transform 1 0 16652 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_181
timestamp 1644511149
transform 1 0 17756 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_193
timestamp 1644511149
transform 1 0 18860 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_205
timestamp 1644511149
transform 1 0 19964 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_217
timestamp 1644511149
transform 1 0 21068 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_223
timestamp 1644511149
transform 1 0 21620 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_225
timestamp 1644511149
transform 1 0 21804 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_237
timestamp 1644511149
transform 1 0 22908 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_249
timestamp 1644511149
transform 1 0 24012 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_261
timestamp 1644511149
transform 1 0 25116 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_273
timestamp 1644511149
transform 1 0 26220 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_279
timestamp 1644511149
transform 1 0 26772 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_281
timestamp 1644511149
transform 1 0 26956 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_293
timestamp 1644511149
transform 1 0 28060 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_305
timestamp 1644511149
transform 1 0 29164 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_317
timestamp 1644511149
transform 1 0 30268 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_329
timestamp 1644511149
transform 1 0 31372 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_335
timestamp 1644511149
transform 1 0 31924 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_337
timestamp 1644511149
transform 1 0 32108 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_349
timestamp 1644511149
transform 1 0 33212 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_361
timestamp 1644511149
transform 1 0 34316 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_373
timestamp 1644511149
transform 1 0 35420 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_377
timestamp 1644511149
transform 1 0 35788 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_115_384
timestamp 1644511149
transform 1 0 36432 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_115_393
timestamp 1644511149
transform 1 0 37260 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_115_401
timestamp 1644511149
transform 1 0 37996 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_405
timestamp 1644511149
transform 1 0 38364 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_417
timestamp 1644511149
transform 1 0 39468 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_429
timestamp 1644511149
transform 1 0 40572 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_441
timestamp 1644511149
transform 1 0 41676 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_447
timestamp 1644511149
transform 1 0 42228 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_449
timestamp 1644511149
transform 1 0 42412 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_461
timestamp 1644511149
transform 1 0 43516 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_473
timestamp 1644511149
transform 1 0 44620 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_485
timestamp 1644511149
transform 1 0 45724 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_497
timestamp 1644511149
transform 1 0 46828 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_503
timestamp 1644511149
transform 1 0 47380 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_505
timestamp 1644511149
transform 1 0 47564 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_517
timestamp 1644511149
transform 1 0 48668 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_529
timestamp 1644511149
transform 1 0 49772 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_541
timestamp 1644511149
transform 1 0 50876 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_553
timestamp 1644511149
transform 1 0 51980 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_559
timestamp 1644511149
transform 1 0 52532 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_561
timestamp 1644511149
transform 1 0 52716 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_573
timestamp 1644511149
transform 1 0 53820 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_585
timestamp 1644511149
transform 1 0 54924 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_597
timestamp 1644511149
transform 1 0 56028 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_609
timestamp 1644511149
transform 1 0 57132 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_615
timestamp 1644511149
transform 1 0 57684 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_617
timestamp 1644511149
transform 1 0 57868 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_629
timestamp 1644511149
transform 1 0 58972 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_641
timestamp 1644511149
transform 1 0 60076 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_653
timestamp 1644511149
transform 1 0 61180 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_665
timestamp 1644511149
transform 1 0 62284 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_671
timestamp 1644511149
transform 1 0 62836 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_673
timestamp 1644511149
transform 1 0 63020 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_685
timestamp 1644511149
transform 1 0 64124 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_697
timestamp 1644511149
transform 1 0 65228 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_709
timestamp 1644511149
transform 1 0 66332 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_721
timestamp 1644511149
transform 1 0 67436 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_727
timestamp 1644511149
transform 1 0 67988 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_115_729
timestamp 1644511149
transform 1 0 68172 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_116_3
timestamp 1644511149
transform 1 0 1380 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_116_7
timestamp 1644511149
transform 1 0 1748 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_14
timestamp 1644511149
transform 1 0 2392 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_24
timestamp 1644511149
transform 1 0 3312 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_116_45
timestamp 1644511149
transform 1 0 5244 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_57
timestamp 1644511149
transform 1 0 6348 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_69
timestamp 1644511149
transform 1 0 7452 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_116_81
timestamp 1644511149
transform 1 0 8556 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_85
timestamp 1644511149
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_97
timestamp 1644511149
transform 1 0 10028 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_109
timestamp 1644511149
transform 1 0 11132 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_121
timestamp 1644511149
transform 1 0 12236 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_133
timestamp 1644511149
transform 1 0 13340 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_139
timestamp 1644511149
transform 1 0 13892 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_141
timestamp 1644511149
transform 1 0 14076 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_153
timestamp 1644511149
transform 1 0 15180 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_165
timestamp 1644511149
transform 1 0 16284 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_177
timestamp 1644511149
transform 1 0 17388 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_189
timestamp 1644511149
transform 1 0 18492 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_195
timestamp 1644511149
transform 1 0 19044 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_197
timestamp 1644511149
transform 1 0 19228 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_209
timestamp 1644511149
transform 1 0 20332 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_221
timestamp 1644511149
transform 1 0 21436 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_233
timestamp 1644511149
transform 1 0 22540 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_245
timestamp 1644511149
transform 1 0 23644 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_251
timestamp 1644511149
transform 1 0 24196 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_253
timestamp 1644511149
transform 1 0 24380 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_265
timestamp 1644511149
transform 1 0 25484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_277
timestamp 1644511149
transform 1 0 26588 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_289
timestamp 1644511149
transform 1 0 27692 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_301
timestamp 1644511149
transform 1 0 28796 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_307
timestamp 1644511149
transform 1 0 29348 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_309
timestamp 1644511149
transform 1 0 29532 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_321
timestamp 1644511149
transform 1 0 30636 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_333
timestamp 1644511149
transform 1 0 31740 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_345
timestamp 1644511149
transform 1 0 32844 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_357
timestamp 1644511149
transform 1 0 33948 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_363
timestamp 1644511149
transform 1 0 34500 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_116_365
timestamp 1644511149
transform 1 0 34684 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_116_369
timestamp 1644511149
transform 1 0 35052 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_386
timestamp 1644511149
transform 1 0 36616 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_398
timestamp 1644511149
transform 1 0 37720 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_410
timestamp 1644511149
transform 1 0 38824 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_116_418
timestamp 1644511149
transform 1 0 39560 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_116_421
timestamp 1644511149
transform 1 0 39836 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_433
timestamp 1644511149
transform 1 0 40940 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_445
timestamp 1644511149
transform 1 0 42044 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_457
timestamp 1644511149
transform 1 0 43148 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_469
timestamp 1644511149
transform 1 0 44252 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_475
timestamp 1644511149
transform 1 0 44804 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_477
timestamp 1644511149
transform 1 0 44988 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_489
timestamp 1644511149
transform 1 0 46092 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_501
timestamp 1644511149
transform 1 0 47196 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_513
timestamp 1644511149
transform 1 0 48300 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_525
timestamp 1644511149
transform 1 0 49404 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_531
timestamp 1644511149
transform 1 0 49956 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_533
timestamp 1644511149
transform 1 0 50140 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_545
timestamp 1644511149
transform 1 0 51244 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_557
timestamp 1644511149
transform 1 0 52348 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_569
timestamp 1644511149
transform 1 0 53452 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_581
timestamp 1644511149
transform 1 0 54556 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_587
timestamp 1644511149
transform 1 0 55108 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_589
timestamp 1644511149
transform 1 0 55292 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_601
timestamp 1644511149
transform 1 0 56396 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_613
timestamp 1644511149
transform 1 0 57500 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_625
timestamp 1644511149
transform 1 0 58604 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_637
timestamp 1644511149
transform 1 0 59708 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_643
timestamp 1644511149
transform 1 0 60260 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_645
timestamp 1644511149
transform 1 0 60444 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_657
timestamp 1644511149
transform 1 0 61548 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_669
timestamp 1644511149
transform 1 0 62652 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_681
timestamp 1644511149
transform 1 0 63756 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_693
timestamp 1644511149
transform 1 0 64860 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_699
timestamp 1644511149
transform 1 0 65412 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_701
timestamp 1644511149
transform 1 0 65596 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_713
timestamp 1644511149
transform 1 0 66700 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_116_717
timestamp 1644511149
transform 1 0 67068 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_116_724
timestamp 1644511149
transform 1 0 67712 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_116_732
timestamp 1644511149
transform 1 0 68448 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_3
timestamp 1644511149
transform 1 0 1380 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_7
timestamp 1644511149
transform 1 0 1748 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_11
timestamp 1644511149
transform 1 0 2116 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_117_31
timestamp 1644511149
transform 1 0 3956 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_117_51
timestamp 1644511149
transform 1 0 5796 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_55
timestamp 1644511149
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_57
timestamp 1644511149
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_69
timestamp 1644511149
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_81
timestamp 1644511149
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_93
timestamp 1644511149
transform 1 0 9660 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_105
timestamp 1644511149
transform 1 0 10764 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_111
timestamp 1644511149
transform 1 0 11316 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_113
timestamp 1644511149
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_125
timestamp 1644511149
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_137
timestamp 1644511149
transform 1 0 13708 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_149
timestamp 1644511149
transform 1 0 14812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_161
timestamp 1644511149
transform 1 0 15916 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_167
timestamp 1644511149
transform 1 0 16468 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_169
timestamp 1644511149
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_181
timestamp 1644511149
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_193
timestamp 1644511149
transform 1 0 18860 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_205
timestamp 1644511149
transform 1 0 19964 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_217
timestamp 1644511149
transform 1 0 21068 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_223
timestamp 1644511149
transform 1 0 21620 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_225
timestamp 1644511149
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_237
timestamp 1644511149
transform 1 0 22908 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_249
timestamp 1644511149
transform 1 0 24012 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_261
timestamp 1644511149
transform 1 0 25116 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_273
timestamp 1644511149
transform 1 0 26220 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_279
timestamp 1644511149
transform 1 0 26772 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_281
timestamp 1644511149
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_293
timestamp 1644511149
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_305
timestamp 1644511149
transform 1 0 29164 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_317
timestamp 1644511149
transform 1 0 30268 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_329
timestamp 1644511149
transform 1 0 31372 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_335
timestamp 1644511149
transform 1 0 31924 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_337
timestamp 1644511149
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_349
timestamp 1644511149
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_361
timestamp 1644511149
transform 1 0 34316 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_373
timestamp 1644511149
transform 1 0 35420 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_377
timestamp 1644511149
transform 1 0 35788 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_384
timestamp 1644511149
transform 1 0 36432 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_393
timestamp 1644511149
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_405
timestamp 1644511149
transform 1 0 38364 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_417
timestamp 1644511149
transform 1 0 39468 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_429
timestamp 1644511149
transform 1 0 40572 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_441
timestamp 1644511149
transform 1 0 41676 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_447
timestamp 1644511149
transform 1 0 42228 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_449
timestamp 1644511149
transform 1 0 42412 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_461
timestamp 1644511149
transform 1 0 43516 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_473
timestamp 1644511149
transform 1 0 44620 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_485
timestamp 1644511149
transform 1 0 45724 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_497
timestamp 1644511149
transform 1 0 46828 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_503
timestamp 1644511149
transform 1 0 47380 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_505
timestamp 1644511149
transform 1 0 47564 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_517
timestamp 1644511149
transform 1 0 48668 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_529
timestamp 1644511149
transform 1 0 49772 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_541
timestamp 1644511149
transform 1 0 50876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_553
timestamp 1644511149
transform 1 0 51980 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_559
timestamp 1644511149
transform 1 0 52532 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_561
timestamp 1644511149
transform 1 0 52716 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_573
timestamp 1644511149
transform 1 0 53820 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_585
timestamp 1644511149
transform 1 0 54924 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_597
timestamp 1644511149
transform 1 0 56028 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_609
timestamp 1644511149
transform 1 0 57132 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_615
timestamp 1644511149
transform 1 0 57684 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_617
timestamp 1644511149
transform 1 0 57868 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_629
timestamp 1644511149
transform 1 0 58972 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_641
timestamp 1644511149
transform 1 0 60076 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_653
timestamp 1644511149
transform 1 0 61180 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_665
timestamp 1644511149
transform 1 0 62284 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_671
timestamp 1644511149
transform 1 0 62836 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_673
timestamp 1644511149
transform 1 0 63020 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_685
timestamp 1644511149
transform 1 0 64124 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_697
timestamp 1644511149
transform 1 0 65228 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_117_724
timestamp 1644511149
transform 1 0 67712 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_117_729
timestamp 1644511149
transform 1 0 68172 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_24
timestamp 1644511149
transform 1 0 3312 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_45
timestamp 1644511149
transform 1 0 5244 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_118_61
timestamp 1644511149
transform 1 0 6716 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_73
timestamp 1644511149
transform 1 0 7820 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_81
timestamp 1644511149
transform 1 0 8556 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_85
timestamp 1644511149
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_97
timestamp 1644511149
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_109
timestamp 1644511149
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_121
timestamp 1644511149
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1644511149
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1644511149
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_141
timestamp 1644511149
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_153
timestamp 1644511149
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_165
timestamp 1644511149
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_177
timestamp 1644511149
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_189
timestamp 1644511149
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_195
timestamp 1644511149
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_197
timestamp 1644511149
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_209
timestamp 1644511149
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_221
timestamp 1644511149
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_233
timestamp 1644511149
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_245
timestamp 1644511149
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_251
timestamp 1644511149
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_253
timestamp 1644511149
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_265
timestamp 1644511149
transform 1 0 25484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_277
timestamp 1644511149
transform 1 0 26588 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_289
timestamp 1644511149
transform 1 0 27692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_301
timestamp 1644511149
transform 1 0 28796 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_307
timestamp 1644511149
transform 1 0 29348 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_309
timestamp 1644511149
transform 1 0 29532 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_321
timestamp 1644511149
transform 1 0 30636 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_333
timestamp 1644511149
transform 1 0 31740 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_345
timestamp 1644511149
transform 1 0 32844 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_357
timestamp 1644511149
transform 1 0 33948 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_363
timestamp 1644511149
transform 1 0 34500 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_365
timestamp 1644511149
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_377
timestamp 1644511149
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_389
timestamp 1644511149
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_401
timestamp 1644511149
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_413
timestamp 1644511149
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_419
timestamp 1644511149
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_421
timestamp 1644511149
transform 1 0 39836 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_433
timestamp 1644511149
transform 1 0 40940 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_445
timestamp 1644511149
transform 1 0 42044 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_457
timestamp 1644511149
transform 1 0 43148 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_469
timestamp 1644511149
transform 1 0 44252 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_475
timestamp 1644511149
transform 1 0 44804 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_477
timestamp 1644511149
transform 1 0 44988 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_489
timestamp 1644511149
transform 1 0 46092 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_501
timestamp 1644511149
transform 1 0 47196 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_513
timestamp 1644511149
transform 1 0 48300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_525
timestamp 1644511149
transform 1 0 49404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_531
timestamp 1644511149
transform 1 0 49956 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_533
timestamp 1644511149
transform 1 0 50140 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_545
timestamp 1644511149
transform 1 0 51244 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_557
timestamp 1644511149
transform 1 0 52348 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_569
timestamp 1644511149
transform 1 0 53452 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_581
timestamp 1644511149
transform 1 0 54556 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_587
timestamp 1644511149
transform 1 0 55108 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_589
timestamp 1644511149
transform 1 0 55292 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_601
timestamp 1644511149
transform 1 0 56396 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_613
timestamp 1644511149
transform 1 0 57500 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_625
timestamp 1644511149
transform 1 0 58604 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_637
timestamp 1644511149
transform 1 0 59708 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_643
timestamp 1644511149
transform 1 0 60260 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_645
timestamp 1644511149
transform 1 0 60444 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_657
timestamp 1644511149
transform 1 0 61548 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_669
timestamp 1644511149
transform 1 0 62652 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_681
timestamp 1644511149
transform 1 0 63756 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_693
timestamp 1644511149
transform 1 0 64860 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_699
timestamp 1644511149
transform 1 0 65412 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_701
timestamp 1644511149
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_713
timestamp 1644511149
transform 1 0 66700 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_118_717
timestamp 1644511149
transform 1 0 67068 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_118_724
timestamp 1644511149
transform 1 0 67712 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_118_732
timestamp 1644511149
transform 1 0 68448 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_119_3
timestamp 1644511149
transform 1 0 1380 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_119_11
timestamp 1644511149
transform 1 0 2116 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_31
timestamp 1644511149
transform 1 0 3956 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_51
timestamp 1644511149
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1644511149
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_57
timestamp 1644511149
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_69
timestamp 1644511149
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_81
timestamp 1644511149
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_93
timestamp 1644511149
transform 1 0 9660 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_105
timestamp 1644511149
transform 1 0 10764 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_111
timestamp 1644511149
transform 1 0 11316 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_113
timestamp 1644511149
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_125
timestamp 1644511149
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_137
timestamp 1644511149
transform 1 0 13708 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_149
timestamp 1644511149
transform 1 0 14812 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_161
timestamp 1644511149
transform 1 0 15916 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_167
timestamp 1644511149
transform 1 0 16468 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_169
timestamp 1644511149
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_181
timestamp 1644511149
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_193
timestamp 1644511149
transform 1 0 18860 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_205
timestamp 1644511149
transform 1 0 19964 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_217
timestamp 1644511149
transform 1 0 21068 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_223
timestamp 1644511149
transform 1 0 21620 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_225
timestamp 1644511149
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_237
timestamp 1644511149
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_249
timestamp 1644511149
transform 1 0 24012 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_261
timestamp 1644511149
transform 1 0 25116 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_273
timestamp 1644511149
transform 1 0 26220 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_279
timestamp 1644511149
transform 1 0 26772 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_281
timestamp 1644511149
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_293
timestamp 1644511149
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_305
timestamp 1644511149
transform 1 0 29164 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_317
timestamp 1644511149
transform 1 0 30268 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_329
timestamp 1644511149
transform 1 0 31372 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_335
timestamp 1644511149
transform 1 0 31924 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_337
timestamp 1644511149
transform 1 0 32108 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_349
timestamp 1644511149
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_361
timestamp 1644511149
transform 1 0 34316 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_373
timestamp 1644511149
transform 1 0 35420 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_385
timestamp 1644511149
transform 1 0 36524 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_391
timestamp 1644511149
transform 1 0 37076 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_393
timestamp 1644511149
transform 1 0 37260 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_405
timestamp 1644511149
transform 1 0 38364 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_417
timestamp 1644511149
transform 1 0 39468 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_429
timestamp 1644511149
transform 1 0 40572 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_441
timestamp 1644511149
transform 1 0 41676 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_447
timestamp 1644511149
transform 1 0 42228 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_449
timestamp 1644511149
transform 1 0 42412 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_461
timestamp 1644511149
transform 1 0 43516 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_473
timestamp 1644511149
transform 1 0 44620 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_485
timestamp 1644511149
transform 1 0 45724 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_497
timestamp 1644511149
transform 1 0 46828 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_503
timestamp 1644511149
transform 1 0 47380 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_505
timestamp 1644511149
transform 1 0 47564 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_517
timestamp 1644511149
transform 1 0 48668 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_529
timestamp 1644511149
transform 1 0 49772 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_541
timestamp 1644511149
transform 1 0 50876 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_553
timestamp 1644511149
transform 1 0 51980 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_559
timestamp 1644511149
transform 1 0 52532 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_561
timestamp 1644511149
transform 1 0 52716 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_573
timestamp 1644511149
transform 1 0 53820 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_585
timestamp 1644511149
transform 1 0 54924 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_597
timestamp 1644511149
transform 1 0 56028 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_609
timestamp 1644511149
transform 1 0 57132 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_615
timestamp 1644511149
transform 1 0 57684 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_617
timestamp 1644511149
transform 1 0 57868 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_629
timestamp 1644511149
transform 1 0 58972 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_641
timestamp 1644511149
transform 1 0 60076 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_653
timestamp 1644511149
transform 1 0 61180 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_665
timestamp 1644511149
transform 1 0 62284 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_671
timestamp 1644511149
transform 1 0 62836 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_673
timestamp 1644511149
transform 1 0 63020 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_685
timestamp 1644511149
transform 1 0 64124 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_697
timestamp 1644511149
transform 1 0 65228 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_119_724
timestamp 1644511149
transform 1 0 67712 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_729
timestamp 1644511149
transform 1 0 68172 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_120_3
timestamp 1644511149
transform 1 0 1380 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_7
timestamp 1644511149
transform 1 0 1748 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_120_24
timestamp 1644511149
transform 1 0 3312 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_120_29
timestamp 1644511149
transform 1 0 3772 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_120_58
timestamp 1644511149
transform 1 0 6440 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_70
timestamp 1644511149
transform 1 0 7544 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_120_82
timestamp 1644511149
transform 1 0 8648 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_120_85
timestamp 1644511149
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_97
timestamp 1644511149
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_109
timestamp 1644511149
transform 1 0 11132 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_121
timestamp 1644511149
transform 1 0 12236 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_133
timestamp 1644511149
transform 1 0 13340 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_139
timestamp 1644511149
transform 1 0 13892 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_141
timestamp 1644511149
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_153
timestamp 1644511149
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_165
timestamp 1644511149
transform 1 0 16284 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_177
timestamp 1644511149
transform 1 0 17388 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_189
timestamp 1644511149
transform 1 0 18492 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_195
timestamp 1644511149
transform 1 0 19044 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_197
timestamp 1644511149
transform 1 0 19228 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_209
timestamp 1644511149
transform 1 0 20332 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_221
timestamp 1644511149
transform 1 0 21436 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_233
timestamp 1644511149
transform 1 0 22540 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_245
timestamp 1644511149
transform 1 0 23644 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_251
timestamp 1644511149
transform 1 0 24196 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_253
timestamp 1644511149
transform 1 0 24380 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_265
timestamp 1644511149
transform 1 0 25484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_277
timestamp 1644511149
transform 1 0 26588 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_289
timestamp 1644511149
transform 1 0 27692 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_301
timestamp 1644511149
transform 1 0 28796 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_307
timestamp 1644511149
transform 1 0 29348 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_309
timestamp 1644511149
transform 1 0 29532 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_321
timestamp 1644511149
transform 1 0 30636 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_333
timestamp 1644511149
transform 1 0 31740 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_345
timestamp 1644511149
transform 1 0 32844 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_357
timestamp 1644511149
transform 1 0 33948 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_363
timestamp 1644511149
transform 1 0 34500 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_365
timestamp 1644511149
transform 1 0 34684 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_377
timestamp 1644511149
transform 1 0 35788 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_389
timestamp 1644511149
transform 1 0 36892 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_120_398
timestamp 1644511149
transform 1 0 37720 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_410
timestamp 1644511149
transform 1 0 38824 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_120_418
timestamp 1644511149
transform 1 0 39560 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_120_421
timestamp 1644511149
transform 1 0 39836 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_120_433
timestamp 1644511149
transform 1 0 40940 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_120_440
timestamp 1644511149
transform 1 0 41584 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_452
timestamp 1644511149
transform 1 0 42688 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_464
timestamp 1644511149
transform 1 0 43792 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_477
timestamp 1644511149
transform 1 0 44988 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_489
timestamp 1644511149
transform 1 0 46092 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_501
timestamp 1644511149
transform 1 0 47196 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_513
timestamp 1644511149
transform 1 0 48300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_525
timestamp 1644511149
transform 1 0 49404 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_531
timestamp 1644511149
transform 1 0 49956 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_536
timestamp 1644511149
transform 1 0 50416 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_548
timestamp 1644511149
transform 1 0 51520 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_560
timestamp 1644511149
transform 1 0 52624 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_572
timestamp 1644511149
transform 1 0 53728 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_120_584
timestamp 1644511149
transform 1 0 54832 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_120_589
timestamp 1644511149
transform 1 0 55292 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_601
timestamp 1644511149
transform 1 0 56396 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_613
timestamp 1644511149
transform 1 0 57500 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_625
timestamp 1644511149
transform 1 0 58604 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_637
timestamp 1644511149
transform 1 0 59708 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_643
timestamp 1644511149
transform 1 0 60260 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_645
timestamp 1644511149
transform 1 0 60444 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_657
timestamp 1644511149
transform 1 0 61548 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_669
timestamp 1644511149
transform 1 0 62652 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_681
timestamp 1644511149
transform 1 0 63756 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_693
timestamp 1644511149
transform 1 0 64860 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_699
timestamp 1644511149
transform 1 0 65412 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_120_701
timestamp 1644511149
transform 1 0 65596 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_120_710
timestamp 1644511149
transform 1 0 66424 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_120_719
timestamp 1644511149
transform 1 0 67252 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_120_729
timestamp 1644511149
transform 1 0 68172 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_121_3
timestamp 1644511149
transform 1 0 1380 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_121_10
timestamp 1644511149
transform 1 0 2024 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_14
timestamp 1644511149
transform 1 0 2392 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_31
timestamp 1644511149
transform 1 0 3956 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_43
timestamp 1644511149
transform 1 0 5060 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1644511149
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_57
timestamp 1644511149
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_69
timestamp 1644511149
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_81
timestamp 1644511149
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_93
timestamp 1644511149
transform 1 0 9660 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_105
timestamp 1644511149
transform 1 0 10764 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_111
timestamp 1644511149
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_113
timestamp 1644511149
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_125
timestamp 1644511149
transform 1 0 12604 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_137
timestamp 1644511149
transform 1 0 13708 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_149
timestamp 1644511149
transform 1 0 14812 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_161
timestamp 1644511149
transform 1 0 15916 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_167
timestamp 1644511149
transform 1 0 16468 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_169
timestamp 1644511149
transform 1 0 16652 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_181
timestamp 1644511149
transform 1 0 17756 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_193
timestamp 1644511149
transform 1 0 18860 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_205
timestamp 1644511149
transform 1 0 19964 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_217
timestamp 1644511149
transform 1 0 21068 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_223
timestamp 1644511149
transform 1 0 21620 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_225
timestamp 1644511149
transform 1 0 21804 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_237
timestamp 1644511149
transform 1 0 22908 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_249
timestamp 1644511149
transform 1 0 24012 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_255
timestamp 1644511149
transform 1 0 24564 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_259
timestamp 1644511149
transform 1 0 24932 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_271
timestamp 1644511149
transform 1 0 26036 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_121_279
timestamp 1644511149
transform 1 0 26772 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_121_281
timestamp 1644511149
transform 1 0 26956 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_121_286
timestamp 1644511149
transform 1 0 27416 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_298
timestamp 1644511149
transform 1 0 28520 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_310
timestamp 1644511149
transform 1 0 29624 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_121_322
timestamp 1644511149
transform 1 0 30728 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_121_328
timestamp 1644511149
transform 1 0 31280 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_121_337
timestamp 1644511149
transform 1 0 32108 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_349
timestamp 1644511149
transform 1 0 33212 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_361
timestamp 1644511149
transform 1 0 34316 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_373
timestamp 1644511149
transform 1 0 35420 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_121_381
timestamp 1644511149
transform 1 0 36156 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_121_387
timestamp 1644511149
transform 1 0 36708 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_391
timestamp 1644511149
transform 1 0 37076 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_121_414
timestamp 1644511149
transform 1 0 39192 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_121_439
timestamp 1644511149
transform 1 0 41492 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_121_447
timestamp 1644511149
transform 1 0 42228 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_121_449
timestamp 1644511149
transform 1 0 42412 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_121_455
timestamp 1644511149
transform 1 0 42964 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_467
timestamp 1644511149
transform 1 0 44068 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_500
timestamp 1644511149
transform 1 0 47104 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_121_505
timestamp 1644511149
transform 1 0 47564 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_517
timestamp 1644511149
transform 1 0 48668 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_121_525
timestamp 1644511149
transform 1 0 49404 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_121_548
timestamp 1644511149
transform 1 0 51520 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_564
timestamp 1644511149
transform 1 0 52992 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_576
timestamp 1644511149
transform 1 0 54096 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_588
timestamp 1644511149
transform 1 0 55200 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_121_596
timestamp 1644511149
transform 1 0 55936 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_121_602
timestamp 1644511149
transform 1 0 56488 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_121_614
timestamp 1644511149
transform 1 0 57592 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_121_638
timestamp 1644511149
transform 1 0 59800 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_650
timestamp 1644511149
transform 1 0 60904 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_656
timestamp 1644511149
transform 1 0 61456 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_660
timestamp 1644511149
transform 1 0 61824 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_673
timestamp 1644511149
transform 1 0 63020 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_685
timestamp 1644511149
transform 1 0 64124 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_121_696
timestamp 1644511149
transform 1 0 65136 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_121_721
timestamp 1644511149
transform 1 0 67436 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_727
timestamp 1644511149
transform 1 0 67988 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_121_729
timestamp 1644511149
transform 1 0 68172 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_122_24
timestamp 1644511149
transform 1 0 3312 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_122_29
timestamp 1644511149
transform 1 0 3772 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_37
timestamp 1644511149
transform 1 0 4508 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_41
timestamp 1644511149
transform 1 0 4876 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_45
timestamp 1644511149
transform 1 0 5244 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_49
timestamp 1644511149
transform 1 0 5612 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_122_74
timestamp 1644511149
transform 1 0 7912 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_122_82
timestamp 1644511149
transform 1 0 8648 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_122_85
timestamp 1644511149
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_97
timestamp 1644511149
transform 1 0 10028 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_122_104
timestamp 1644511149
transform 1 0 10672 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_122_129
timestamp 1644511149
transform 1 0 12972 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_137
timestamp 1644511149
transform 1 0 13708 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_122_141
timestamp 1644511149
transform 1 0 14076 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_122_153
timestamp 1644511149
transform 1 0 15180 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_159
timestamp 1644511149
transform 1 0 15732 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_122_184
timestamp 1644511149
transform 1 0 18032 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_197
timestamp 1644511149
transform 1 0 19228 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_209
timestamp 1644511149
transform 1 0 20332 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_221
timestamp 1644511149
transform 1 0 21436 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_233
timestamp 1644511149
transform 1 0 22540 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_245
timestamp 1644511149
transform 1 0 23644 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_251
timestamp 1644511149
transform 1 0 24196 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_122_253
timestamp 1644511149
transform 1 0 24380 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_277
timestamp 1644511149
transform 1 0 26588 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_281
timestamp 1644511149
transform 1 0 26956 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_303
timestamp 1644511149
transform 1 0 28980 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_307
timestamp 1644511149
transform 1 0 29348 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_309
timestamp 1644511149
transform 1 0 29532 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_321
timestamp 1644511149
transform 1 0 30636 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_122_346
timestamp 1644511149
transform 1 0 32936 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_358
timestamp 1644511149
transform 1 0 34040 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_122_365
timestamp 1644511149
transform 1 0 34684 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_377
timestamp 1644511149
transform 1 0 35788 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_381
timestamp 1644511149
transform 1 0 36156 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_403
timestamp 1644511149
transform 1 0 38180 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_122_414
timestamp 1644511149
transform 1 0 39192 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_122_421
timestamp 1644511149
transform 1 0 39836 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_425
timestamp 1644511149
transform 1 0 40204 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_447
timestamp 1644511149
transform 1 0 42228 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_122_472
timestamp 1644511149
transform 1 0 44528 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_122_477
timestamp 1644511149
transform 1 0 44988 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_122_483
timestamp 1644511149
transform 1 0 45540 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_491
timestamp 1644511149
transform 1 0 46276 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_513
timestamp 1644511149
transform 1 0 48300 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_517
timestamp 1644511149
transform 1 0 48668 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_521
timestamp 1644511149
transform 1 0 49036 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_122_528
timestamp 1644511149
transform 1 0 49680 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_122_533
timestamp 1644511149
transform 1 0 50140 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_557
timestamp 1644511149
transform 1 0 52348 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_122_582
timestamp 1644511149
transform 1 0 54648 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_122_589
timestamp 1644511149
transform 1 0 55292 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_122_597
timestamp 1644511149
transform 1 0 56028 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_122_620
timestamp 1644511149
transform 1 0 58144 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_632
timestamp 1644511149
transform 1 0 59248 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_636
timestamp 1644511149
transform 1 0 59616 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_640
timestamp 1644511149
transform 1 0 59984 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_122_666
timestamp 1644511149
transform 1 0 62376 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_122_691
timestamp 1644511149
transform 1 0 64676 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_699
timestamp 1644511149
transform 1 0 65412 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_704
timestamp 1644511149
transform 1 0 65872 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_122_729
timestamp 1644511149
transform 1 0 68172 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_9
timestamp 1644511149
transform 1 0 1932 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_123_16
timestamp 1644511149
transform 1 0 2576 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_29
timestamp 1644511149
transform 1 0 3772 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_123_37
timestamp 1644511149
transform 1 0 4508 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_41
timestamp 1644511149
transform 1 0 4876 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_53
timestamp 1644511149
transform 1 0 5980 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_60
timestamp 1644511149
transform 1 0 6624 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_123_72
timestamp 1644511149
transform 1 0 7728 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_123_77
timestamp 1644511149
transform 1 0 8188 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_83
timestamp 1644511149
transform 1 0 8740 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_85
timestamp 1644511149
transform 1 0 8924 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_97
timestamp 1644511149
transform 1 0 10028 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_109
timestamp 1644511149
transform 1 0 11132 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_116
timestamp 1644511149
transform 1 0 11776 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_128
timestamp 1644511149
transform 1 0 12880 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_141
timestamp 1644511149
transform 1 0 14076 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_123_149
timestamp 1644511149
transform 1 0 14812 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_161
timestamp 1644511149
transform 1 0 15916 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_167
timestamp 1644511149
transform 1 0 16468 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_172
timestamp 1644511149
transform 1 0 16928 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_184
timestamp 1644511149
transform 1 0 18032 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_197
timestamp 1644511149
transform 1 0 19228 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_123_205
timestamp 1644511149
transform 1 0 19964 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_123_217
timestamp 1644511149
transform 1 0 21068 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_223
timestamp 1644511149
transform 1 0 21620 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_225
timestamp 1644511149
transform 1 0 21804 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_237
timestamp 1644511149
transform 1 0 22908 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_249
timestamp 1644511149
transform 1 0 24012 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_123_253
timestamp 1644511149
transform 1 0 24380 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_259
timestamp 1644511149
transform 1 0 24932 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_271
timestamp 1644511149
transform 1 0 26036 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_123_279
timestamp 1644511149
transform 1 0 26772 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_123_281
timestamp 1644511149
transform 1 0 26956 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_123_286
timestamp 1644511149
transform 1 0 27416 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_298
timestamp 1644511149
transform 1 0 28520 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_123_306
timestamp 1644511149
transform 1 0 29256 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_123_309
timestamp 1644511149
transform 1 0 29532 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_321
timestamp 1644511149
transform 1 0 30636 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_123_328
timestamp 1644511149
transform 1 0 31280 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_123_337
timestamp 1644511149
transform 1 0 32108 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_349
timestamp 1644511149
transform 1 0 33212 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_361
timestamp 1644511149
transform 1 0 34316 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_123_365
timestamp 1644511149
transform 1 0 34684 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_123_373
timestamp 1644511149
transform 1 0 35420 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_123_380
timestamp 1644511149
transform 1 0 36064 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_387
timestamp 1644511149
transform 1 0 36708 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_391
timestamp 1644511149
transform 1 0 37076 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_123_393
timestamp 1644511149
transform 1 0 37260 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_397
timestamp 1644511149
transform 1 0 37628 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_123_409
timestamp 1644511149
transform 1 0 38732 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_123_413
timestamp 1644511149
transform 1 0 39100 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_419
timestamp 1644511149
transform 1 0 39652 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_421
timestamp 1644511149
transform 1 0 39836 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_433
timestamp 1644511149
transform 1 0 40940 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_123_439
timestamp 1644511149
transform 1 0 41492 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_123_447
timestamp 1644511149
transform 1 0 42228 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_123_449
timestamp 1644511149
transform 1 0 42412 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_455
timestamp 1644511149
transform 1 0 42964 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_467
timestamp 1644511149
transform 1 0 44068 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_123_475
timestamp 1644511149
transform 1 0 44804 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_123_477
timestamp 1644511149
transform 1 0 44988 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_123_483
timestamp 1644511149
transform 1 0 45540 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_490
timestamp 1644511149
transform 1 0 46184 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_123_497
timestamp 1644511149
transform 1 0 46828 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_503
timestamp 1644511149
transform 1 0 47380 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_505
timestamp 1644511149
transform 1 0 47564 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_517
timestamp 1644511149
transform 1 0 48668 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_529
timestamp 1644511149
transform 1 0 49772 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_123_533
timestamp 1644511149
transform 1 0 50140 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_123_540
timestamp 1644511149
transform 1 0 50784 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_552
timestamp 1644511149
transform 1 0 51888 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_123_564
timestamp 1644511149
transform 1 0 52992 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_576
timestamp 1644511149
transform 1 0 54096 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_589
timestamp 1644511149
transform 1 0 55292 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_123_595
timestamp 1644511149
transform 1 0 55844 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_599
timestamp 1644511149
transform 1 0 56212 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_123_603
timestamp 1644511149
transform 1 0 56580 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_123_612
timestamp 1644511149
transform 1 0 57408 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_123_620
timestamp 1644511149
transform 1 0 58144 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_632
timestamp 1644511149
transform 1 0 59248 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_648
timestamp 1644511149
transform 1 0 60720 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_660
timestamp 1644511149
transform 1 0 61824 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_123_665
timestamp 1644511149
transform 1 0 62284 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_671
timestamp 1644511149
transform 1 0 62836 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_673
timestamp 1644511149
transform 1 0 63020 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_123_685
timestamp 1644511149
transform 1 0 64124 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_123_689
timestamp 1644511149
transform 1 0 64492 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_696
timestamp 1644511149
transform 1 0 65136 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_123_701
timestamp 1644511149
transform 1 0 65596 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_123_724
timestamp 1644511149
transform 1 0 67712 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_729
timestamp 1644511149
transform 1 0 68172 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 68816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 68816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 68816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 68816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 68816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 68816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 68816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 68816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 68816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 68816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 68816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 68816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 68816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 68816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 68816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 68816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 68816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 68816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 68816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 68816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 68816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 68816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 68816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 68816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 68816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 68816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 68816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 68816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 68816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 68816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 68816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 68816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 68816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 68816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 68816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 68816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 68816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 68816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 68816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 68816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 68816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 68816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 68816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 68816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 68816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 68816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 68816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 68816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 68816 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 68816 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 68816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 68816 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 68816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 68816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 68816 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 68816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 68816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 68816 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 68816 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 68816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 68816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 68816 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 68816 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 68816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 68816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 68816 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 68816 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 68816 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 68816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 68816 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 68816 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 68816 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 68816 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 68816 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 68816 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 68816 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 68816 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 68816 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 68816 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 68816 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 68816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 68816 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 68816 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1644511149
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1644511149
transform -1 0 68816 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1644511149
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1644511149
transform -1 0 68816 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1644511149
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1644511149
transform -1 0 68816 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1644511149
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1644511149
transform -1 0 68816 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1644511149
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1644511149
transform -1 0 68816 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1644511149
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1644511149
transform -1 0 68816 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1644511149
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1644511149
transform -1 0 68816 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1644511149
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1644511149
transform -1 0 68816 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1644511149
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1644511149
transform -1 0 68816 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1644511149
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1644511149
transform -1 0 68816 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1644511149
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1644511149
transform -1 0 68816 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1644511149
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1644511149
transform -1 0 68816 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1644511149
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1644511149
transform -1 0 68816 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1644511149
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1644511149
transform -1 0 68816 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1644511149
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1644511149
transform -1 0 68816 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1644511149
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1644511149
transform -1 0 68816 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1644511149
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1644511149
transform -1 0 68816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1644511149
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1644511149
transform -1 0 68816 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1644511149
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1644511149
transform -1 0 68816 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1644511149
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1644511149
transform -1 0 68816 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1644511149
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1644511149
transform -1 0 68816 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1644511149
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1644511149
transform -1 0 68816 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1644511149
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1644511149
transform -1 0 68816 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1644511149
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1644511149
transform -1 0 68816 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1644511149
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1644511149
transform -1 0 68816 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1644511149
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1644511149
transform -1 0 68816 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1644511149
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1644511149
transform -1 0 68816 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1644511149
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1644511149
transform -1 0 68816 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1644511149
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1644511149
transform -1 0 68816 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1644511149
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1644511149
transform -1 0 68816 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1644511149
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1644511149
transform -1 0 68816 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1644511149
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1644511149
transform -1 0 68816 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1644511149
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1644511149
transform -1 0 68816 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1644511149
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1644511149
transform -1 0 68816 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1644511149
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1644511149
transform -1 0 68816 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1644511149
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1644511149
transform -1 0 68816 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1644511149
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1644511149
transform -1 0 68816 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1644511149
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1644511149
transform -1 0 68816 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1644511149
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1644511149
transform -1 0 68816 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1644511149
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1644511149
transform -1 0 68816 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1644511149
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1644511149
transform -1 0 68816 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1644511149
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1644511149
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1644511149
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1644511149
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1644511149
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1644511149
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1644511149
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1644511149
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1644511149
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1644511149
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1644511149
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1644511149
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1644511149
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1644511149
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1644511149
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1644511149
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1644511149
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1644511149
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1644511149
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1644511149
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1644511149
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1644511149
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1644511149
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1644511149
transform 1 0 62928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1644511149
transform 1 0 68080 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1644511149
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1644511149
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1644511149
transform 1 0 60352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1644511149
transform 1 0 65504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1644511149
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1644511149
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1644511149
transform 1 0 62928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1644511149
transform 1 0 68080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1644511149
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1644511149
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1644511149
transform 1 0 60352 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1644511149
transform 1 0 65504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1644511149
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1644511149
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1644511149
transform 1 0 62928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1644511149
transform 1 0 68080 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1644511149
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1644511149
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1644511149
transform 1 0 60352 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1644511149
transform 1 0 65504 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1644511149
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1644511149
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1644511149
transform 1 0 62928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1644511149
transform 1 0 68080 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1644511149
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1644511149
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1644511149
transform 1 0 60352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1644511149
transform 1 0 65504 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1644511149
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1644511149
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1644511149
transform 1 0 62928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1644511149
transform 1 0 68080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1644511149
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1644511149
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1644511149
transform 1 0 60352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1644511149
transform 1 0 65504 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1644511149
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1644511149
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1644511149
transform 1 0 62928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1644511149
transform 1 0 68080 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1644511149
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1644511149
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1644511149
transform 1 0 60352 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1644511149
transform 1 0 65504 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1644511149
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1644511149
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1644511149
transform 1 0 62928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1644511149
transform 1 0 68080 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1644511149
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1644511149
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1644511149
transform 1 0 60352 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1644511149
transform 1 0 65504 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1644511149
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1644511149
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1644511149
transform 1 0 62928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1644511149
transform 1 0 68080 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1644511149
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1644511149
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1644511149
transform 1 0 60352 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1644511149
transform 1 0 65504 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1644511149
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1644511149
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1644511149
transform 1 0 62928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1644511149
transform 1 0 68080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1644511149
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1644511149
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1644511149
transform 1 0 60352 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1644511149
transform 1 0 65504 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1644511149
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1644511149
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1644511149
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1644511149
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1644511149
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1644511149
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1644511149
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1644511149
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1644511149
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1644511149
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1644511149
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1644511149
transform 1 0 62928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1644511149
transform 1 0 68080 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1644511149
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1644511149
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1644511149
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1644511149
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1644511149
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1644511149
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1644511149
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1644511149
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1644511149
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1644511149
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1644511149
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1644511149
transform 1 0 60352 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1644511149
transform 1 0 65504 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1644511149
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1644511149
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1644511149
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1644511149
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1644511149
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1644511149
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1644511149
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1644511149
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1644511149
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1644511149
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1644511149
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1644511149
transform 1 0 62928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1644511149
transform 1 0 68080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1644511149
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1644511149
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1644511149
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1644511149
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1644511149
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1644511149
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1644511149
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1644511149
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1644511149
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1644511149
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1644511149
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1644511149
transform 1 0 60352 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1644511149
transform 1 0 65504 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1644511149
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1644511149
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1644511149
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1644511149
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1644511149
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1644511149
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1644511149
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1644511149
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1644511149
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1644511149
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1644511149
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1644511149
transform 1 0 62928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1644511149
transform 1 0 68080 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1644511149
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1644511149
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1644511149
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1644511149
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1644511149
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1644511149
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1644511149
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1644511149
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1644511149
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1644511149
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1644511149
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1644511149
transform 1 0 60352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1644511149
transform 1 0 65504 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1644511149
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1644511149
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1644511149
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1644511149
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1644511149
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1644511149
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1644511149
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1644511149
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1644511149
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1644511149
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1644511149
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1644511149
transform 1 0 62928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1644511149
transform 1 0 68080 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1644511149
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1644511149
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1644511149
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1644511149
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1644511149
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1644511149
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1644511149
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1644511149
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1644511149
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1644511149
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1644511149
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1644511149
transform 1 0 60352 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1644511149
transform 1 0 65504 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1644511149
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1644511149
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1644511149
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1644511149
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1644511149
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1644511149
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1644511149
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1644511149
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1644511149
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1644511149
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1644511149
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1644511149
transform 1 0 62928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1644511149
transform 1 0 68080 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1644511149
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1644511149
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1644511149
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1644511149
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1644511149
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1644511149
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1644511149
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1644511149
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1644511149
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1644511149
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1644511149
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1644511149
transform 1 0 60352 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1644511149
transform 1 0 65504 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1644511149
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1644511149
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1644511149
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1644511149
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1644511149
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1644511149
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1644511149
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1644511149
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1644511149
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1644511149
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1644511149
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1644511149
transform 1 0 62928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1644511149
transform 1 0 68080 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1644511149
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1644511149
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1644511149
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1644511149
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1644511149
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1644511149
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1644511149
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1644511149
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1644511149
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1644511149
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1644511149
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1644511149
transform 1 0 60352 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1644511149
transform 1 0 65504 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1644511149
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1644511149
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1644511149
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1644511149
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1644511149
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1644511149
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1644511149
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1644511149
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1644511149
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1644511149
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1644511149
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1644511149
transform 1 0 62928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1644511149
transform 1 0 68080 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1644511149
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1644511149
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1644511149
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1644511149
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1644511149
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1644511149
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1644511149
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1644511149
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1644511149
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1644511149
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1644511149
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1644511149
transform 1 0 60352 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1644511149
transform 1 0 65504 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1644511149
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1644511149
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1644511149
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1644511149
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1644511149
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1644511149
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1644511149
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1644511149
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1644511149
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1644511149
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1644511149
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1644511149
transform 1 0 62928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1644511149
transform 1 0 68080 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1644511149
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1644511149
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1644511149
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1644511149
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1644511149
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1644511149
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1644511149
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1644511149
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1644511149
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1644511149
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1644511149
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1644511149
transform 1 0 60352 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1644511149
transform 1 0 65504 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1644511149
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1644511149
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1644511149
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1644511149
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1644511149
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1644511149
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1644511149
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1644511149
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1644511149
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1644511149
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1644511149
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1644511149
transform 1 0 62928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1644511149
transform 1 0 68080 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1644511149
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1644511149
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1644511149
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1644511149
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1644511149
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1644511149
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1644511149
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1644511149
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1644511149
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1644511149
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1644511149
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1644511149
transform 1 0 60352 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1644511149
transform 1 0 65504 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1644511149
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1644511149
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1644511149
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1644511149
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1644511149
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1644511149
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1644511149
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1644511149
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1644511149
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1644511149
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1644511149
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1644511149
transform 1 0 62928 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1644511149
transform 1 0 68080 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1644511149
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1644511149
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1644511149
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1644511149
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1644511149
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1644511149
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1644511149
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1644511149
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1644511149
transform 1 0 44896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1644511149
transform 1 0 50048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1644511149
transform 1 0 55200 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1644511149
transform 1 0 60352 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1644511149
transform 1 0 65504 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1644511149
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1644511149
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1644511149
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1644511149
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1644511149
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1644511149
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1644511149
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1644511149
transform 1 0 42320 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1644511149
transform 1 0 47472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1644511149
transform 1 0 52624 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1644511149
transform 1 0 57776 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1644511149
transform 1 0 62928 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1644511149
transform 1 0 68080 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1644511149
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1644511149
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1644511149
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1644511149
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1644511149
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1644511149
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1644511149
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1644511149
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1644511149
transform 1 0 44896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1644511149
transform 1 0 50048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1644511149
transform 1 0 55200 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1644511149
transform 1 0 60352 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1644511149
transform 1 0 65504 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1644511149
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1644511149
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1644511149
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1644511149
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1644511149
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1644511149
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1644511149
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1644511149
transform 1 0 42320 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1644511149
transform 1 0 47472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1644511149
transform 1 0 52624 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1644511149
transform 1 0 57776 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1637
timestamp 1644511149
transform 1 0 62928 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1638
timestamp 1644511149
transform 1 0 68080 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1639
timestamp 1644511149
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1640
timestamp 1644511149
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1641
timestamp 1644511149
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1642
timestamp 1644511149
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1643
timestamp 1644511149
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1644
timestamp 1644511149
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1645
timestamp 1644511149
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1646
timestamp 1644511149
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1647
timestamp 1644511149
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1648
timestamp 1644511149
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1649
timestamp 1644511149
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1650
timestamp 1644511149
transform 1 0 60352 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1651
timestamp 1644511149
transform 1 0 65504 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1652
timestamp 1644511149
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1653
timestamp 1644511149
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1654
timestamp 1644511149
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1655
timestamp 1644511149
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1656
timestamp 1644511149
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1657
timestamp 1644511149
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1658
timestamp 1644511149
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1659
timestamp 1644511149
transform 1 0 42320 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1660
timestamp 1644511149
transform 1 0 47472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1661
timestamp 1644511149
transform 1 0 52624 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1662
timestamp 1644511149
transform 1 0 57776 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1663
timestamp 1644511149
transform 1 0 62928 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1664
timestamp 1644511149
transform 1 0 68080 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1665
timestamp 1644511149
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1666
timestamp 1644511149
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1667
timestamp 1644511149
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1668
timestamp 1644511149
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1669
timestamp 1644511149
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1670
timestamp 1644511149
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1671
timestamp 1644511149
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1672
timestamp 1644511149
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1673
timestamp 1644511149
transform 1 0 44896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1674
timestamp 1644511149
transform 1 0 50048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1675
timestamp 1644511149
transform 1 0 55200 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1676
timestamp 1644511149
transform 1 0 60352 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1677
timestamp 1644511149
transform 1 0 65504 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1678
timestamp 1644511149
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1679
timestamp 1644511149
transform 1 0 11408 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1680
timestamp 1644511149
transform 1 0 16560 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1681
timestamp 1644511149
transform 1 0 21712 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1682
timestamp 1644511149
transform 1 0 26864 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1683
timestamp 1644511149
transform 1 0 32016 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1684
timestamp 1644511149
transform 1 0 37168 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1685
timestamp 1644511149
transform 1 0 42320 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1686
timestamp 1644511149
transform 1 0 47472 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1687
timestamp 1644511149
transform 1 0 52624 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1688
timestamp 1644511149
transform 1 0 57776 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1689
timestamp 1644511149
transform 1 0 62928 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1690
timestamp 1644511149
transform 1 0 68080 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1691
timestamp 1644511149
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1692
timestamp 1644511149
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1693
timestamp 1644511149
transform 1 0 13984 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1694
timestamp 1644511149
transform 1 0 19136 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1695
timestamp 1644511149
transform 1 0 24288 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1696
timestamp 1644511149
transform 1 0 29440 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1697
timestamp 1644511149
transform 1 0 34592 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1698
timestamp 1644511149
transform 1 0 39744 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1699
timestamp 1644511149
transform 1 0 44896 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1700
timestamp 1644511149
transform 1 0 50048 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1701
timestamp 1644511149
transform 1 0 55200 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1702
timestamp 1644511149
transform 1 0 60352 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1703
timestamp 1644511149
transform 1 0 65504 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1704
timestamp 1644511149
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1705
timestamp 1644511149
transform 1 0 11408 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1706
timestamp 1644511149
transform 1 0 16560 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1707
timestamp 1644511149
transform 1 0 21712 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1708
timestamp 1644511149
transform 1 0 26864 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1709
timestamp 1644511149
transform 1 0 32016 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1710
timestamp 1644511149
transform 1 0 37168 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1711
timestamp 1644511149
transform 1 0 42320 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1712
timestamp 1644511149
transform 1 0 47472 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1713
timestamp 1644511149
transform 1 0 52624 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1714
timestamp 1644511149
transform 1 0 57776 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1715
timestamp 1644511149
transform 1 0 62928 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1716
timestamp 1644511149
transform 1 0 68080 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1717
timestamp 1644511149
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1718
timestamp 1644511149
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1719
timestamp 1644511149
transform 1 0 13984 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1720
timestamp 1644511149
transform 1 0 19136 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1721
timestamp 1644511149
transform 1 0 24288 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1722
timestamp 1644511149
transform 1 0 29440 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1723
timestamp 1644511149
transform 1 0 34592 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1724
timestamp 1644511149
transform 1 0 39744 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1725
timestamp 1644511149
transform 1 0 44896 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1726
timestamp 1644511149
transform 1 0 50048 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1727
timestamp 1644511149
transform 1 0 55200 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1728
timestamp 1644511149
transform 1 0 60352 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1729
timestamp 1644511149
transform 1 0 65504 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1730
timestamp 1644511149
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1731
timestamp 1644511149
transform 1 0 11408 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1732
timestamp 1644511149
transform 1 0 16560 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1733
timestamp 1644511149
transform 1 0 21712 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1734
timestamp 1644511149
transform 1 0 26864 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1735
timestamp 1644511149
transform 1 0 32016 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1736
timestamp 1644511149
transform 1 0 37168 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1737
timestamp 1644511149
transform 1 0 42320 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1738
timestamp 1644511149
transform 1 0 47472 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1739
timestamp 1644511149
transform 1 0 52624 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1740
timestamp 1644511149
transform 1 0 57776 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1741
timestamp 1644511149
transform 1 0 62928 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1742
timestamp 1644511149
transform 1 0 68080 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1743
timestamp 1644511149
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1744
timestamp 1644511149
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1745
timestamp 1644511149
transform 1 0 13984 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1746
timestamp 1644511149
transform 1 0 19136 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1747
timestamp 1644511149
transform 1 0 24288 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1748
timestamp 1644511149
transform 1 0 29440 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1749
timestamp 1644511149
transform 1 0 34592 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1750
timestamp 1644511149
transform 1 0 39744 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1751
timestamp 1644511149
transform 1 0 44896 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1752
timestamp 1644511149
transform 1 0 50048 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1753
timestamp 1644511149
transform 1 0 55200 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1754
timestamp 1644511149
transform 1 0 60352 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1755
timestamp 1644511149
transform 1 0 65504 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1756
timestamp 1644511149
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1757
timestamp 1644511149
transform 1 0 11408 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1758
timestamp 1644511149
transform 1 0 16560 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1759
timestamp 1644511149
transform 1 0 21712 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1760
timestamp 1644511149
transform 1 0 26864 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1761
timestamp 1644511149
transform 1 0 32016 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1762
timestamp 1644511149
transform 1 0 37168 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1763
timestamp 1644511149
transform 1 0 42320 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1764
timestamp 1644511149
transform 1 0 47472 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1765
timestamp 1644511149
transform 1 0 52624 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1766
timestamp 1644511149
transform 1 0 57776 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1767
timestamp 1644511149
transform 1 0 62928 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1768
timestamp 1644511149
transform 1 0 68080 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1769
timestamp 1644511149
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1770
timestamp 1644511149
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1771
timestamp 1644511149
transform 1 0 13984 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1772
timestamp 1644511149
transform 1 0 19136 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1773
timestamp 1644511149
transform 1 0 24288 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1774
timestamp 1644511149
transform 1 0 29440 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1775
timestamp 1644511149
transform 1 0 34592 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1776
timestamp 1644511149
transform 1 0 39744 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1777
timestamp 1644511149
transform 1 0 44896 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1778
timestamp 1644511149
transform 1 0 50048 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1779
timestamp 1644511149
transform 1 0 55200 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1780
timestamp 1644511149
transform 1 0 60352 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1781
timestamp 1644511149
transform 1 0 65504 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1782
timestamp 1644511149
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1783
timestamp 1644511149
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1784
timestamp 1644511149
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1785
timestamp 1644511149
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1786
timestamp 1644511149
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1787
timestamp 1644511149
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1788
timestamp 1644511149
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1789
timestamp 1644511149
transform 1 0 42320 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1790
timestamp 1644511149
transform 1 0 47472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1791
timestamp 1644511149
transform 1 0 52624 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1792
timestamp 1644511149
transform 1 0 57776 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1793
timestamp 1644511149
transform 1 0 62928 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1794
timestamp 1644511149
transform 1 0 68080 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1795
timestamp 1644511149
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1796
timestamp 1644511149
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1797
timestamp 1644511149
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1798
timestamp 1644511149
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1799
timestamp 1644511149
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1800
timestamp 1644511149
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1801
timestamp 1644511149
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1802
timestamp 1644511149
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1803
timestamp 1644511149
transform 1 0 44896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1804
timestamp 1644511149
transform 1 0 50048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1805
timestamp 1644511149
transform 1 0 55200 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1806
timestamp 1644511149
transform 1 0 60352 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1807
timestamp 1644511149
transform 1 0 65504 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1808
timestamp 1644511149
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1809
timestamp 1644511149
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1810
timestamp 1644511149
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1811
timestamp 1644511149
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1812
timestamp 1644511149
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1813
timestamp 1644511149
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1814
timestamp 1644511149
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1815
timestamp 1644511149
transform 1 0 42320 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1816
timestamp 1644511149
transform 1 0 47472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1817
timestamp 1644511149
transform 1 0 52624 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1818
timestamp 1644511149
transform 1 0 57776 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1819
timestamp 1644511149
transform 1 0 62928 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1820
timestamp 1644511149
transform 1 0 68080 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1821
timestamp 1644511149
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1822
timestamp 1644511149
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1823
timestamp 1644511149
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1824
timestamp 1644511149
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1825
timestamp 1644511149
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1826
timestamp 1644511149
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1827
timestamp 1644511149
transform 1 0 34592 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1828
timestamp 1644511149
transform 1 0 39744 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1829
timestamp 1644511149
transform 1 0 44896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1830
timestamp 1644511149
transform 1 0 50048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1831
timestamp 1644511149
transform 1 0 55200 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1832
timestamp 1644511149
transform 1 0 60352 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1833
timestamp 1644511149
transform 1 0 65504 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1834
timestamp 1644511149
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1835
timestamp 1644511149
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1836
timestamp 1644511149
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1837
timestamp 1644511149
transform 1 0 21712 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1838
timestamp 1644511149
transform 1 0 26864 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1839
timestamp 1644511149
transform 1 0 32016 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1840
timestamp 1644511149
transform 1 0 37168 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1841
timestamp 1644511149
transform 1 0 42320 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1842
timestamp 1644511149
transform 1 0 47472 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1843
timestamp 1644511149
transform 1 0 52624 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1844
timestamp 1644511149
transform 1 0 57776 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1845
timestamp 1644511149
transform 1 0 62928 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1846
timestamp 1644511149
transform 1 0 68080 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1847
timestamp 1644511149
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1848
timestamp 1644511149
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1849
timestamp 1644511149
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1850
timestamp 1644511149
transform 1 0 19136 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1851
timestamp 1644511149
transform 1 0 24288 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1852
timestamp 1644511149
transform 1 0 29440 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1853
timestamp 1644511149
transform 1 0 34592 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1854
timestamp 1644511149
transform 1 0 39744 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1855
timestamp 1644511149
transform 1 0 44896 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1856
timestamp 1644511149
transform 1 0 50048 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1857
timestamp 1644511149
transform 1 0 55200 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1858
timestamp 1644511149
transform 1 0 60352 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1859
timestamp 1644511149
transform 1 0 65504 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1860
timestamp 1644511149
transform 1 0 3680 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1861
timestamp 1644511149
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1862
timestamp 1644511149
transform 1 0 8832 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1863
timestamp 1644511149
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1864
timestamp 1644511149
transform 1 0 13984 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1865
timestamp 1644511149
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1866
timestamp 1644511149
transform 1 0 19136 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1867
timestamp 1644511149
transform 1 0 21712 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1868
timestamp 1644511149
transform 1 0 24288 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1869
timestamp 1644511149
transform 1 0 26864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1870
timestamp 1644511149
transform 1 0 29440 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1871
timestamp 1644511149
transform 1 0 32016 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1872
timestamp 1644511149
transform 1 0 34592 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1873
timestamp 1644511149
transform 1 0 37168 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1874
timestamp 1644511149
transform 1 0 39744 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1875
timestamp 1644511149
transform 1 0 42320 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1876
timestamp 1644511149
transform 1 0 44896 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1877
timestamp 1644511149
transform 1 0 47472 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1878
timestamp 1644511149
transform 1 0 50048 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1879
timestamp 1644511149
transform 1 0 52624 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1880
timestamp 1644511149
transform 1 0 55200 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1881
timestamp 1644511149
transform 1 0 57776 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1882
timestamp 1644511149
transform 1 0 60352 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1883
timestamp 1644511149
transform 1 0 62928 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1884
timestamp 1644511149
transform 1 0 65504 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1885
timestamp 1644511149
transform 1 0 68080 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1179_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23552 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1180_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38548 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1181_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38272 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1182_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39928 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1183_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42872 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1184_
timestamp 1644511149
transform 1 0 43240 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1185_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42412 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_2  _1186_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42228 0 1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _1187_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43148 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1188_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44896 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1189_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43516 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _1190_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42780 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1191_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41308 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1192_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41400 0 1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1193_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41032 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1194_
timestamp 1644511149
transform 1 0 41216 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1195_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42964 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1196_
timestamp 1644511149
transform 1 0 42964 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1197_
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1198_
timestamp 1644511149
transform 1 0 43516 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1199_
timestamp 1644511149
transform 1 0 44160 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1200_
timestamp 1644511149
transform 1 0 43424 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1201_
timestamp 1644511149
transform 1 0 43424 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1202_
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1203_
timestamp 1644511149
transform 1 0 40480 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1204_
timestamp 1644511149
transform 1 0 41492 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1205_
timestamp 1644511149
transform 1 0 42780 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1206_
timestamp 1644511149
transform 1 0 41584 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1207_
timestamp 1644511149
transform 1 0 43332 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1208_
timestamp 1644511149
transform 1 0 43976 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1209_
timestamp 1644511149
transform 1 0 42780 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1210_
timestamp 1644511149
transform 1 0 43700 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1211_
timestamp 1644511149
transform 1 0 43792 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1212_
timestamp 1644511149
transform 1 0 44436 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1213_
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1214_
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1215_
timestamp 1644511149
transform 1 0 40112 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1216_
timestamp 1644511149
transform 1 0 40388 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1217_
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1218_
timestamp 1644511149
transform 1 0 38732 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1219_
timestamp 1644511149
transform 1 0 38180 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1220_
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1221_
timestamp 1644511149
transform 1 0 39652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1222_
timestamp 1644511149
transform 1 0 38916 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1223_
timestamp 1644511149
transform 1 0 38272 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1224_
timestamp 1644511149
transform 1 0 39100 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1225_
timestamp 1644511149
transform 1 0 38916 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1226_
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1227_
timestamp 1644511149
transform 1 0 39560 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1228_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1229_
timestamp 1644511149
transform 1 0 43884 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1230_
timestamp 1644511149
transform 1 0 44160 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1231_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41400 0 1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1232_
timestamp 1644511149
transform 1 0 40572 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_4  _1233_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38732 0 -1 47872
box -38 -48 1602 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1234_
timestamp 1644511149
transform 1 0 29348 0 -1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1235_
timestamp 1644511149
transform 1 0 29716 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1236_
timestamp 1644511149
transform 1 0 31096 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1237_
timestamp 1644511149
transform 1 0 27600 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1238_
timestamp 1644511149
transform 1 0 26956 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1239_
timestamp 1644511149
transform 1 0 27140 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1240_
timestamp 1644511149
transform 1 0 26496 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1241_
timestamp 1644511149
transform 1 0 27416 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1242_
timestamp 1644511149
transform 1 0 27140 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1243_
timestamp 1644511149
transform 1 0 27232 0 -1 60928
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1244_
timestamp 1644511149
transform 1 0 26220 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1245_
timestamp 1644511149
transform 1 0 15916 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1246_
timestamp 1644511149
transform 1 0 22172 0 -1 60928
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1247_
timestamp 1644511149
transform 1 0 22172 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1248_
timestamp 1644511149
transform 1 0 14720 0 -1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1249_
timestamp 1644511149
transform 1 0 14444 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1250_
timestamp 1644511149
transform 1 0 14996 0 1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1251_
timestamp 1644511149
transform 1 0 14904 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1252_
timestamp 1644511149
transform 1 0 14904 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1253_
timestamp 1644511149
transform 1 0 14628 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1254_
timestamp 1644511149
transform 1 0 14444 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1255_
timestamp 1644511149
transform 1 0 14076 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1256_
timestamp 1644511149
transform 1 0 14996 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1257_
timestamp 1644511149
transform 1 0 14996 0 1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1258_
timestamp 1644511149
transform 1 0 14352 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1259_
timestamp 1644511149
transform 1 0 14904 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1260_
timestamp 1644511149
transform 1 0 14996 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1261_
timestamp 1644511149
transform 1 0 15088 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1262_
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1263_
timestamp 1644511149
transform 1 0 15272 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1264_
timestamp 1644511149
transform 1 0 15180 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1265_
timestamp 1644511149
transform 1 0 15364 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1266_
timestamp 1644511149
transform 1 0 15456 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1267_
timestamp 1644511149
transform 1 0 23092 0 1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1268_
timestamp 1644511149
transform 1 0 23092 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1269_
timestamp 1644511149
transform 1 0 42412 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _1270_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42964 0 1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1271_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43700 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1272_
timestamp 1644511149
transform 1 0 45724 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1273_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45448 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1274_
timestamp 1644511149
transform 1 0 45448 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1275_
timestamp 1644511149
transform 1 0 38180 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1276_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42872 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1277_
timestamp 1644511149
transform 1 0 27968 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1278_
timestamp 1644511149
transform 1 0 28060 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1279_
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1280_
timestamp 1644511149
transform 1 0 28336 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1281_
timestamp 1644511149
transform 1 0 28888 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1282_
timestamp 1644511149
transform 1 0 29808 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1283_
timestamp 1644511149
transform 1 0 30636 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1284_
timestamp 1644511149
transform 1 0 29624 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1285_
timestamp 1644511149
transform 1 0 30452 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1286_
timestamp 1644511149
transform 1 0 28060 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1287_
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1288_
timestamp 1644511149
transform 1 0 34040 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1289_
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1290_
timestamp 1644511149
transform 1 0 34040 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1291_
timestamp 1644511149
transform 1 0 33764 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1292_
timestamp 1644511149
transform 1 0 35420 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1293_
timestamp 1644511149
transform 1 0 32936 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1294_
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1295_
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1296_
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1297_
timestamp 1644511149
transform 1 0 32476 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1298_
timestamp 1644511149
transform 1 0 32200 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1299_
timestamp 1644511149
transform 1 0 24472 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1300_
timestamp 1644511149
transform 1 0 22632 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1301_
timestamp 1644511149
transform 1 0 22264 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1302_
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1303_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1304_
timestamp 1644511149
transform 1 0 23000 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1305_
timestamp 1644511149
transform 1 0 22816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1306_
timestamp 1644511149
transform 1 0 23092 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1307_
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1308_
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1309_
timestamp 1644511149
transform 1 0 23000 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1310_
timestamp 1644511149
transform 1 0 26956 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1311_
timestamp 1644511149
transform 1 0 26036 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1312_
timestamp 1644511149
transform 1 0 50232 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1313_
timestamp 1644511149
transform 1 0 50324 0 1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1314_
timestamp 1644511149
transform 1 0 48668 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1315_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47748 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1316_
timestamp 1644511149
transform 1 0 50140 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1317_
timestamp 1644511149
transform 1 0 43700 0 -1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_2  _1318_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 48024 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__or4b_1  _1319_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1320_
timestamp 1644511149
transform 1 0 44252 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1321_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44528 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1322_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39284 0 -1 50048
box -38 -48 1234 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1323_
timestamp 1644511149
transform 1 0 25116 0 -1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1324_
timestamp 1644511149
transform 1 0 25300 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1325_
timestamp 1644511149
transform 1 0 25208 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1326_
timestamp 1644511149
transform 1 0 25300 0 -1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1327_
timestamp 1644511149
transform 1 0 25208 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1328_
timestamp 1644511149
transform 1 0 25024 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1329_
timestamp 1644511149
transform 1 0 25300 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1330_
timestamp 1644511149
transform 1 0 25208 0 -1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1331_
timestamp 1644511149
transform 1 0 25208 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1332_
timestamp 1644511149
transform 1 0 25116 0 -1 59840
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1333_
timestamp 1644511149
transform 1 0 24932 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1334_
timestamp 1644511149
transform 1 0 16652 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1335_
timestamp 1644511149
transform 1 0 17388 0 1 59840
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1336_
timestamp 1644511149
transform 1 0 17388 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1337_
timestamp 1644511149
transform 1 0 16652 0 -1 59840
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1338_
timestamp 1644511149
transform 1 0 15916 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1339_
timestamp 1644511149
transform 1 0 17020 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1340_
timestamp 1644511149
transform 1 0 16928 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1341_
timestamp 1644511149
transform 1 0 15732 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1342_
timestamp 1644511149
transform 1 0 16652 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1343_
timestamp 1644511149
transform 1 0 15640 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1344_
timestamp 1644511149
transform 1 0 14996 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1345_
timestamp 1644511149
transform 1 0 17020 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1346_
timestamp 1644511149
transform 1 0 13064 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1347_
timestamp 1644511149
transform 1 0 12972 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1348_
timestamp 1644511149
transform 1 0 12972 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1349_
timestamp 1644511149
transform 1 0 12696 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1350_
timestamp 1644511149
transform 1 0 13156 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1351_
timestamp 1644511149
transform 1 0 12972 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1352_
timestamp 1644511149
transform 1 0 13156 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1353_
timestamp 1644511149
transform 1 0 13156 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1354_
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1355_
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1356_
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1357_
timestamp 1644511149
transform 1 0 23644 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1358_
timestamp 1644511149
transform 1 0 50048 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1359_
timestamp 1644511149
transform 1 0 49312 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1360_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1361_
timestamp 1644511149
transform 1 0 44988 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1362_
timestamp 1644511149
transform 1 0 39836 0 1 48960
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _1363_
timestamp 1644511149
transform 1 0 26128 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1364_
timestamp 1644511149
transform 1 0 25300 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1365_
timestamp 1644511149
transform 1 0 25024 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1366_
timestamp 1644511149
transform 1 0 24840 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1367_
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1368_
timestamp 1644511149
transform 1 0 25024 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1369_
timestamp 1644511149
transform 1 0 24748 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1370_
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1371_
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1372_
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1374_
timestamp 1644511149
transform 1 0 30728 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1375_
timestamp 1644511149
transform 1 0 31188 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1376_
timestamp 1644511149
transform 1 0 31280 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1377_
timestamp 1644511149
transform 1 0 31096 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1378_
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1379_
timestamp 1644511149
transform 1 0 31004 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1380_
timestamp 1644511149
transform 1 0 30912 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1381_
timestamp 1644511149
transform 1 0 31556 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1382_
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1383_
timestamp 1644511149
transform 1 0 31188 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1384_
timestamp 1644511149
transform 1 0 31188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1385_
timestamp 1644511149
transform 1 0 25576 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1386_
timestamp 1644511149
transform 1 0 25484 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1387_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1388_
timestamp 1644511149
transform 1 0 25300 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1389_
timestamp 1644511149
transform 1 0 25208 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1390_
timestamp 1644511149
transform 1 0 25300 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1391_
timestamp 1644511149
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1392_
timestamp 1644511149
transform 1 0 24472 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1393_
timestamp 1644511149
transform 1 0 24656 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1394_
timestamp 1644511149
transform 1 0 24472 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1395_
timestamp 1644511149
transform 1 0 24656 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1396_
timestamp 1644511149
transform 1 0 27140 0 -1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1397_
timestamp 1644511149
transform 1 0 27140 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1398_
timestamp 1644511149
transform 1 0 47564 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1399_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43516 0 -1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1400_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 48484 0 -1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1401_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47012 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1402_
timestamp 1644511149
transform 1 0 43240 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1403_
timestamp 1644511149
transform 1 0 44896 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1404_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43332 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1405_
timestamp 1644511149
transform 1 0 27968 0 1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1406_
timestamp 1644511149
transform 1 0 27968 0 -1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1407_
timestamp 1644511149
transform 1 0 27600 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1408_
timestamp 1644511149
transform 1 0 28612 0 1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1409_
timestamp 1644511149
transform 1 0 27416 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1410_
timestamp 1644511149
transform 1 0 28428 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1411_
timestamp 1644511149
transform 1 0 28520 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1412_
timestamp 1644511149
transform 1 0 28244 0 1 60928
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1413_
timestamp 1644511149
transform 1 0 28796 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1414_
timestamp 1644511149
transform 1 0 27324 0 1 60928
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1415_
timestamp 1644511149
transform 1 0 26404 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1416_
timestamp 1644511149
transform 1 0 20424 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1417_
timestamp 1644511149
transform 1 0 20332 0 1 60928
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1418_
timestamp 1644511149
transform 1 0 21068 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1419_
timestamp 1644511149
transform 1 0 19412 0 1 60928
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1420_
timestamp 1644511149
transform 1 0 19504 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1421_
timestamp 1644511149
transform 1 0 18032 0 1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1422_
timestamp 1644511149
transform 1 0 16928 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1423_
timestamp 1644511149
transform 1 0 18768 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1424_
timestamp 1644511149
transform 1 0 17664 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1425_
timestamp 1644511149
transform 1 0 17940 0 1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1426_
timestamp 1644511149
transform 1 0 17388 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1427_
timestamp 1644511149
transform 1 0 19872 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1428_
timestamp 1644511149
transform 1 0 18124 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1429_
timestamp 1644511149
transform 1 0 16836 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1430_
timestamp 1644511149
transform 1 0 17020 0 -1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1431_
timestamp 1644511149
transform 1 0 17020 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1432_
timestamp 1644511149
transform 1 0 17296 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1433_
timestamp 1644511149
transform 1 0 18308 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1434_
timestamp 1644511149
transform 1 0 17572 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1435_
timestamp 1644511149
transform 1 0 17388 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1436_
timestamp 1644511149
transform 1 0 19504 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1437_
timestamp 1644511149
transform 1 0 19412 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1438_
timestamp 1644511149
transform 1 0 24564 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1439_
timestamp 1644511149
transform 1 0 25392 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1440_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35052 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1441_
timestamp 1644511149
transform 1 0 34132 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1442_
timestamp 1644511149
transform 1 0 45356 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1443_
timestamp 1644511149
transform 1 0 48760 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1444_
timestamp 1644511149
transform 1 0 45356 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1445_
timestamp 1644511149
transform 1 0 47564 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a2111oi_1  _1446_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 48300 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1447_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1448_
timestamp 1644511149
transform 1 0 46000 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1449_
timestamp 1644511149
transform 1 0 44804 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_2  _1450_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45632 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1451_
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1452_
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1453_
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1454_
timestamp 1644511149
transform 1 0 30728 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1455_
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1456_
timestamp 1644511149
transform 1 0 32384 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1458_
timestamp 1644511149
transform 1 0 33764 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1459_
timestamp 1644511149
transform 1 0 33764 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1460_
timestamp 1644511149
transform 1 0 33764 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1462_
timestamp 1644511149
transform 1 0 33212 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1463_
timestamp 1644511149
transform 1 0 32844 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1464_
timestamp 1644511149
transform 1 0 32568 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1465_
timestamp 1644511149
transform 1 0 33120 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1466_
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1467_
timestamp 1644511149
transform 1 0 33028 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1468_
timestamp 1644511149
transform 1 0 33120 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1469_
timestamp 1644511149
transform 1 0 32936 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1470_
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1471_
timestamp 1644511149
transform 1 0 33212 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1472_
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1473_
timestamp 1644511149
transform 1 0 32568 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1474_
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1475_
timestamp 1644511149
transform 1 0 27232 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1476_
timestamp 1644511149
transform 1 0 28520 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1477_
timestamp 1644511149
transform 1 0 27784 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1478_
timestamp 1644511149
transform 1 0 28336 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1479_
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1480_
timestamp 1644511149
transform 1 0 26496 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1481_
timestamp 1644511149
transform 1 0 28060 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1482_
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1483_
timestamp 1644511149
transform 1 0 27048 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1484_
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1485_
timestamp 1644511149
transform 1 0 27140 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1486_
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1487_
timestamp 1644511149
transform 1 0 29900 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1488_
timestamp 1644511149
transform 1 0 29072 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1489_
timestamp 1644511149
transform 1 0 28612 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1490_
timestamp 1644511149
transform 1 0 46276 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1491_
timestamp 1644511149
transform 1 0 45908 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1492_
timestamp 1644511149
transform 1 0 46184 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1493_
timestamp 1644511149
transform 1 0 46092 0 -1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1494_
timestamp 1644511149
transform 1 0 30636 0 -1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1495_
timestamp 1644511149
transform 1 0 32108 0 -1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1644511149
transform 1 0 30912 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1497_
timestamp 1644511149
transform 1 0 29808 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1498_
timestamp 1644511149
transform 1 0 30636 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1499_
timestamp 1644511149
transform 1 0 30360 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 1644511149
transform 1 0 31372 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1501_
timestamp 1644511149
transform 1 0 29900 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1502_
timestamp 1644511149
transform 1 0 31096 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1503_
timestamp 1644511149
transform 1 0 20884 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1504_
timestamp 1644511149
transform 1 0 29532 0 1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1505_
timestamp 1644511149
transform 1 0 29532 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1506_
timestamp 1644511149
transform 1 0 21528 0 1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1507_
timestamp 1644511149
transform 1 0 20884 0 -1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1508_
timestamp 1644511149
transform 1 0 21436 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1509_
timestamp 1644511149
transform 1 0 19780 0 1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1510_
timestamp 1644511149
transform 1 0 19964 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1511_
timestamp 1644511149
transform 1 0 19872 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1512_
timestamp 1644511149
transform 1 0 20332 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1513_
timestamp 1644511149
transform 1 0 19780 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1514_
timestamp 1644511149
transform 1 0 20148 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1515_
timestamp 1644511149
transform 1 0 21068 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1516_
timestamp 1644511149
transform 1 0 19688 0 -1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1517_
timestamp 1644511149
transform 1 0 19688 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1518_
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1519_
timestamp 1644511149
transform 1 0 19872 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1520_
timestamp 1644511149
transform 1 0 19504 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1521_
timestamp 1644511149
transform 1 0 19596 0 1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1522_
timestamp 1644511149
transform 1 0 19596 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1523_
timestamp 1644511149
transform 1 0 19688 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1524_
timestamp 1644511149
transform 1 0 20792 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1525_
timestamp 1644511149
transform 1 0 20516 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1526_
timestamp 1644511149
transform 1 0 19964 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1527_
timestamp 1644511149
transform 1 0 37444 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1528_
timestamp 1644511149
transform 1 0 32752 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1529_
timestamp 1644511149
transform 1 0 21896 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1530_
timestamp 1644511149
transform 1 0 22540 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1531_
timestamp 1644511149
transform 1 0 25576 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1532_
timestamp 1644511149
transform 1 0 25760 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1533_
timestamp 1644511149
transform 1 0 45264 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1534_
timestamp 1644511149
transform 1 0 46092 0 1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1535_
timestamp 1644511149
transform 1 0 46092 0 1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _1536_
timestamp 1644511149
transform 1 0 45632 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1537_
timestamp 1644511149
transform 1 0 30176 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1538_
timestamp 1644511149
transform 1 0 29440 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1539_
timestamp 1644511149
transform 1 0 28336 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1540_
timestamp 1644511149
transform 1 0 30360 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1541_
timestamp 1644511149
transform 1 0 30728 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1542_
timestamp 1644511149
transform 1 0 32660 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1543_
timestamp 1644511149
transform 1 0 33856 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1544_
timestamp 1644511149
transform 1 0 35328 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1545_
timestamp 1644511149
transform 1 0 35144 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1546_
timestamp 1644511149
transform 1 0 35236 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1547_
timestamp 1644511149
transform 1 0 35144 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1548_
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1549_
timestamp 1644511149
transform 1 0 35420 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1550_
timestamp 1644511149
transform 1 0 36156 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1551_
timestamp 1644511149
transform 1 0 36340 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1552_
timestamp 1644511149
transform 1 0 35604 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1553_
timestamp 1644511149
transform 1 0 34960 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1554_
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1644511149
transform 1 0 36432 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1556_
timestamp 1644511149
transform 1 0 35696 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1557_
timestamp 1644511149
transform 1 0 35328 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1558_
timestamp 1644511149
transform 1 0 35328 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1559_
timestamp 1644511149
transform 1 0 35052 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1560_
timestamp 1644511149
transform 1 0 35880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1561_
timestamp 1644511149
transform 1 0 29716 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1562_
timestamp 1644511149
transform 1 0 28796 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1563_
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1564_
timestamp 1644511149
transform 1 0 27968 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1565_
timestamp 1644511149
transform 1 0 27508 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1566_
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1567_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1568_
timestamp 1644511149
transform 1 0 33488 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1569_
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1570_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1571_
timestamp 1644511149
transform 1 0 29808 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1572_
timestamp 1644511149
transform 1 0 29624 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1573_
timestamp 1644511149
transform 1 0 30176 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1574_
timestamp 1644511149
transform 1 0 31096 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1575_
timestamp 1644511149
transform 1 0 36064 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _1576_
timestamp 1644511149
transform 1 0 37628 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1577_
timestamp 1644511149
transform 1 0 39928 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1578_
timestamp 1644511149
transform 1 0 40756 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1579_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41216 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1580_
timestamp 1644511149
transform 1 0 36340 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1581_
timestamp 1644511149
transform 1 0 38916 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1582_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41032 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1583_
timestamp 1644511149
transform 1 0 41584 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1584_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42412 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1585_
timestamp 1644511149
transform 1 0 40480 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _1586_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41308 0 -1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1587_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43700 0 1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1588_
timestamp 1644511149
transform 1 0 43608 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1589_
timestamp 1644511149
transform 1 0 44988 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1590_
timestamp 1644511149
transform 1 0 45816 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1591_
timestamp 1644511149
transform 1 0 48760 0 1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1592_
timestamp 1644511149
transform 1 0 48116 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1593_
timestamp 1644511149
transform 1 0 47564 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1594_
timestamp 1644511149
transform 1 0 50140 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1595_
timestamp 1644511149
transform 1 0 50140 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1596_
timestamp 1644511149
transform 1 0 48576 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1597_
timestamp 1644511149
transform 1 0 48300 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1598_
timestamp 1644511149
transform 1 0 49864 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1599_
timestamp 1644511149
transform 1 0 51060 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1600_
timestamp 1644511149
transform 1 0 49864 0 -1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1601_
timestamp 1644511149
transform 1 0 50692 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1602_
timestamp 1644511149
transform 1 0 45448 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1603_
timestamp 1644511149
transform 1 0 45632 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1604_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46092 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1605_
timestamp 1644511149
transform 1 0 37628 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1606_
timestamp 1644511149
transform 1 0 43976 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1607_
timestamp 1644511149
transform 1 0 45816 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1608_
timestamp 1644511149
transform 1 0 49864 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1609_
timestamp 1644511149
transform 1 0 50232 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1610_
timestamp 1644511149
transform 1 0 51060 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1611_
timestamp 1644511149
transform 1 0 51244 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1612_
timestamp 1644511149
transform 1 0 52716 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1613_
timestamp 1644511149
transform 1 0 50876 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1614_
timestamp 1644511149
transform 1 0 51888 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1615_
timestamp 1644511149
transform 1 0 50600 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1616_
timestamp 1644511149
transform 1 0 51428 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1617_
timestamp 1644511149
transform 1 0 51520 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1618_
timestamp 1644511149
transform 1 0 51428 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1619_
timestamp 1644511149
transform 1 0 48852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1620_
timestamp 1644511149
transform 1 0 49220 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1621_
timestamp 1644511149
transform 1 0 47564 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1622_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 48300 0 -1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1623_
timestamp 1644511149
transform 1 0 48300 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1624_
timestamp 1644511149
transform 1 0 46736 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1625_
timestamp 1644511149
transform 1 0 37076 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1626_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46920 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1627_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1628_
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1629_
timestamp 1644511149
transform 1 0 47932 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1630_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1631_
timestamp 1644511149
transform 1 0 48300 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1632_
timestamp 1644511149
transform 1 0 45540 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1633_
timestamp 1644511149
transform 1 0 46368 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1634_
timestamp 1644511149
transform 1 0 43976 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1635_
timestamp 1644511149
transform 1 0 43792 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1636_
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1637_
timestamp 1644511149
transform 1 0 39836 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1638_
timestamp 1644511149
transform 1 0 40664 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1639_
timestamp 1644511149
transform 1 0 39376 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1640_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40664 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1641_
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1642_
timestamp 1644511149
transform 1 0 39836 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1643_
timestamp 1644511149
transform 1 0 41400 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1644_
timestamp 1644511149
transform 1 0 23276 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  _1645_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  _1646_
timestamp 1644511149
transform 1 0 25024 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1647_
timestamp 1644511149
transform 1 0 24288 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1648_
timestamp 1644511149
transform 1 0 33028 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1649_
timestamp 1644511149
transform 1 0 29716 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1650_
timestamp 1644511149
transform 1 0 33580 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1651_
timestamp 1644511149
transform 1 0 33672 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1652_
timestamp 1644511149
transform 1 0 5428 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1653_
timestamp 1644511149
transform 1 0 5980 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1654_
timestamp 1644511149
transform 1 0 66332 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1655_
timestamp 1644511149
transform 1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1656_
timestamp 1644511149
transform 1 0 67160 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1657_
timestamp 1644511149
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1658_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1564 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  _1659_
timestamp 1644511149
transform 1 0 2484 0 -1 67456
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1660_
timestamp 1644511149
transform 1 0 1748 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1661_
timestamp 1644511149
transform 1 0 36432 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1662_
timestamp 1644511149
transform 1 0 67436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1663_
timestamp 1644511149
transform 1 0 67528 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1664_
timestamp 1644511149
transform 1 0 1748 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1665_
timestamp 1644511149
transform 1 0 2484 0 -1 68544
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1666_
timestamp 1644511149
transform 1 0 67252 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1667_
timestamp 1644511149
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1668_
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1669_
timestamp 1644511149
transform 1 0 1932 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1670_
timestamp 1644511149
transform 1 0 42688 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1671_
timestamp 1644511149
transform 1 0 1840 0 1 67456
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1672_
timestamp 1644511149
transform 1 0 66976 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1673_
timestamp 1644511149
transform 1 0 2300 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1674_
timestamp 1644511149
transform 1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1675_
timestamp 1644511149
transform 1 0 24656 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1676_
timestamp 1644511149
transform 1 0 67528 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1677_
timestamp 1644511149
transform 1 0 2484 0 -1 66368
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1678_
timestamp 1644511149
transform 1 0 59708 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1679_
timestamp 1644511149
transform 1 0 2208 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1680_
timestamp 1644511149
transform 1 0 60720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1681_
timestamp 1644511149
transform 1 0 65596 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1682_
timestamp 1644511149
transform 1 0 46552 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1683_
timestamp 1644511149
transform 1 0 4324 0 -1 67456
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1684_
timestamp 1644511149
transform 1 0 67436 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1685_
timestamp 1644511149
transform 1 0 2300 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1686_
timestamp 1644511149
transform 1 0 67436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1687_
timestamp 1644511149
transform 1 0 67528 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1688_
timestamp 1644511149
transform 1 0 41308 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1689_
timestamp 1644511149
transform 1 0 2760 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1690_
timestamp 1644511149
transform 1 0 4048 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1691_
timestamp 1644511149
transform 1 0 49404 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1692_
timestamp 1644511149
transform 1 0 2116 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1644511149
transform 1 0 45264 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1694_
timestamp 1644511149
transform 1 0 15456 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1695_
timestamp 1644511149
transform 1 0 27140 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1696_
timestamp 1644511149
transform 1 0 3772 0 1 66368
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1697_
timestamp 1644511149
transform 1 0 37444 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1698_
timestamp 1644511149
transform 1 0 67344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1699_
timestamp 1644511149
transform 1 0 2760 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1700_
timestamp 1644511149
transform 1 0 67528 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1701_
timestamp 1644511149
transform 1 0 66884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1702_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5612 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1703_
timestamp 1644511149
transform 1 0 1932 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1704_
timestamp 1644511149
transform 1 0 10396 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1705_
timestamp 1644511149
transform 1 0 67160 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1706_
timestamp 1644511149
transform 1 0 1932 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1707_
timestamp 1644511149
transform 1 0 5336 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1708_
timestamp 1644511149
transform 1 0 3772 0 1 65280
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1709_
timestamp 1644511149
transform 1 0 67436 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1710_
timestamp 1644511149
transform 1 0 67436 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1711_
timestamp 1644511149
transform 1 0 2668 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1712_
timestamp 1644511149
transform 1 0 50140 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1713_
timestamp 1644511149
transform 1 0 61916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1714_
timestamp 1644511149
transform 1 0 4324 0 -1 66368
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1715_
timestamp 1644511149
transform 1 0 52716 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1716_
timestamp 1644511149
transform 1 0 67436 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1717_
timestamp 1644511149
transform 1 0 67436 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1718_
timestamp 1644511149
transform 1 0 67528 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1719_
timestamp 1644511149
transform 1 0 2576 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1720_
timestamp 1644511149
transform 1 0 23000 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  _1721_
timestamp 1644511149
transform 1 0 24380 0 1 62016
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1722_
timestamp 1644511149
transform 1 0 33396 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1723_
timestamp 1644511149
transform 1 0 61548 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1724_
timestamp 1644511149
transform 1 0 2024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1725_
timestamp 1644511149
transform 1 0 2392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1726_
timestamp 1644511149
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1727_
timestamp 1644511149
transform 1 0 23920 0 -1 63104
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1728_
timestamp 1644511149
transform 1 0 67436 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1729_
timestamp 1644511149
transform 1 0 56212 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1730_
timestamp 1644511149
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1731_
timestamp 1644511149
transform 1 0 21988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1732_
timestamp 1644511149
transform 1 0 67436 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1733_
timestamp 1644511149
transform 1 0 22448 0 1 62016
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1734_
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1735_
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1736_
timestamp 1644511149
transform 1 0 31004 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1737_
timestamp 1644511149
transform 1 0 4600 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1738_
timestamp 1644511149
transform 1 0 66148 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1739_
timestamp 1644511149
transform 1 0 24380 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1740_
timestamp 1644511149
transform 1 0 38916 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1741_
timestamp 1644511149
transform 1 0 67528 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1742_
timestamp 1644511149
transform 1 0 67436 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1743_
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1744_
timestamp 1644511149
transform 1 0 57868 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1745_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1746_
timestamp 1644511149
transform 1 0 67252 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1747_
timestamp 1644511149
transform 1 0 50140 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1748_
timestamp 1644511149
transform 1 0 32568 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1749_
timestamp 1644511149
transform 1 0 28428 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1750_
timestamp 1644511149
transform 1 0 23460 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1751_
timestamp 1644511149
transform 1 0 23184 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1752_
timestamp 1644511149
transform 1 0 22632 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1753_
timestamp 1644511149
transform 1 0 19780 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1754_
timestamp 1644511149
transform 1 0 23552 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1755_
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1756_
timestamp 1644511149
transform 1 0 19596 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1757_
timestamp 1644511149
transform 1 0 45448 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1758_
timestamp 1644511149
transform 1 0 48668 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1759_
timestamp 1644511149
transform 1 0 48760 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1760_
timestamp 1644511149
transform 1 0 49312 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1761_
timestamp 1644511149
transform 1 0 48760 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1762_
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1763_
timestamp 1644511149
transform 1 0 44988 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1764_
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1765_
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1766_
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1767_
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1768_
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1769_
timestamp 1644511149
transform 1 0 23276 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1770_
timestamp 1644511149
transform 1 0 40204 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1771_
timestamp 1644511149
transform 1 0 24380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1772_
timestamp 1644511149
transform 1 0 23092 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1773_
timestamp 1644511149
transform 1 0 40848 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1774_
timestamp 1644511149
transform 1 0 22632 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1775_
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1776_
timestamp 1644511149
transform 1 0 1840 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1777_
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1778_
timestamp 1644511149
transform 1 0 38824 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1779_
timestamp 1644511149
transform 1 0 38548 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1780_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36892 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1781_
timestamp 1644511149
transform 1 0 17296 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1782_
timestamp 1644511149
transform 1 0 25852 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1783_
timestamp 1644511149
transform 1 0 26128 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _1784_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _1785_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  _1786_
timestamp 1644511149
transform 1 0 36248 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1787_
timestamp 1644511149
transform 1 0 20700 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _1788_
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1789_
timestamp 1644511149
transform 1 0 20516 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _1790_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18952 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _1791_
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  _1792_
timestamp 1644511149
transform 1 0 36616 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1793_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37904 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _1794_
timestamp 1644511149
transform 1 0 38640 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1795_
timestamp 1644511149
transform 1 0 38272 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1796_
timestamp 1644511149
transform 1 0 42412 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1797_
timestamp 1644511149
transform 1 0 38732 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1798_
timestamp 1644511149
transform 1 0 40480 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _1799_
timestamp 1644511149
transform 1 0 42504 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1800_
timestamp 1644511149
transform 1 0 43332 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1801_
timestamp 1644511149
transform 1 0 44988 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1802_
timestamp 1644511149
transform 1 0 36524 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1803_
timestamp 1644511149
transform 1 0 36156 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1804_
timestamp 1644511149
transform 1 0 36708 0 1 63104
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1805_
timestamp 1644511149
transform 1 0 36156 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1806_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36064 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1807_
timestamp 1644511149
transform 1 0 35328 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1808_
timestamp 1644511149
transform 1 0 37260 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1809_
timestamp 1644511149
transform 1 0 36340 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1810_
timestamp 1644511149
transform 1 0 35696 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1811_
timestamp 1644511149
transform 1 0 35696 0 -1 60928
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1812_
timestamp 1644511149
transform 1 0 35236 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1813_
timestamp 1644511149
transform 1 0 34776 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1814_
timestamp 1644511149
transform 1 0 35328 0 -1 63104
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1815_
timestamp 1644511149
transform 1 0 35788 0 -1 62016
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1816_
timestamp 1644511149
transform 1 0 35604 0 1 63104
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1817_
timestamp 1644511149
transform 1 0 34684 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1818_
timestamp 1644511149
transform 1 0 37628 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1819_
timestamp 1644511149
transform 1 0 37720 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1820_
timestamp 1644511149
transform 1 0 36340 0 -1 64192
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1821_
timestamp 1644511149
transform 1 0 37536 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1822_
timestamp 1644511149
transform 1 0 36892 0 1 64192
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1823_
timestamp 1644511149
transform 1 0 38088 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1824_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35880 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1825_
timestamp 1644511149
transform 1 0 35880 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1826_
timestamp 1644511149
transform 1 0 32292 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1827_
timestamp 1644511149
transform 1 0 38548 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1828_
timestamp 1644511149
transform 1 0 36432 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1829_
timestamp 1644511149
transform 1 0 28704 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1830_
timestamp 1644511149
transform 1 0 28428 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1831_
timestamp 1644511149
transform 1 0 36064 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_4  _1832_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37352 0 1 46784
box -38 -48 1786 592
use sky130_fd_sc_hd__o2111a_1  _1833_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35328 0 -1 53312
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1834_
timestamp 1644511149
transform 1 0 36524 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _1835_
timestamp 1644511149
transform 1 0 35696 0 1 55488
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1836_
timestamp 1644511149
transform 1 0 35512 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1837_
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1838_
timestamp 1644511149
transform 1 0 33580 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1839_
timestamp 1644511149
transform 1 0 32844 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1840_
timestamp 1644511149
transform 1 0 29992 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1841_
timestamp 1644511149
transform 1 0 28704 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1842_
timestamp 1644511149
transform 1 0 19044 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1843_
timestamp 1644511149
transform 1 0 33764 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1844_
timestamp 1644511149
transform 1 0 34592 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1845_
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1846_
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1847_
timestamp 1644511149
transform 1 0 36800 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1848_
timestamp 1644511149
transform 1 0 36432 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1849_
timestamp 1644511149
transform 1 0 36248 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1850_
timestamp 1644511149
transform 1 0 38088 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1851_
timestamp 1644511149
transform 1 0 37444 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1852_
timestamp 1644511149
transform 1 0 36984 0 1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1853_
timestamp 1644511149
transform 1 0 36524 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1854_
timestamp 1644511149
transform 1 0 35788 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1855_
timestamp 1644511149
transform 1 0 35512 0 -1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1856_
timestamp 1644511149
transform 1 0 35236 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1857_
timestamp 1644511149
transform 1 0 34224 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1858_
timestamp 1644511149
transform 1 0 34592 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1859_
timestamp 1644511149
transform 1 0 35420 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1860_
timestamp 1644511149
transform 1 0 34132 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1861_
timestamp 1644511149
transform 1 0 34684 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1862_
timestamp 1644511149
transform 1 0 35604 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1863_
timestamp 1644511149
transform 1 0 34684 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1864_
timestamp 1644511149
transform 1 0 35144 0 -1 52224
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1865_
timestamp 1644511149
transform 1 0 35052 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1866_
timestamp 1644511149
transform 1 0 35052 0 1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1867_
timestamp 1644511149
transform 1 0 33580 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1868_
timestamp 1644511149
transform 1 0 37260 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1869_
timestamp 1644511149
transform 1 0 35972 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1870_
timestamp 1644511149
transform 1 0 33948 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1871_
timestamp 1644511149
transform 1 0 39376 0 -1 59840
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_1  _1872_
timestamp 1644511149
transform 1 0 38548 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1873_
timestamp 1644511149
transform 1 0 38548 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1874_
timestamp 1644511149
transform 1 0 39744 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1875_
timestamp 1644511149
transform 1 0 38732 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1876_
timestamp 1644511149
transform 1 0 39836 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1877_
timestamp 1644511149
transform 1 0 39836 0 1 58752
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1878_
timestamp 1644511149
transform 1 0 39928 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1879_
timestamp 1644511149
transform 1 0 38640 0 1 58752
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1880_
timestamp 1644511149
transform 1 0 37168 0 1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1881_
timestamp 1644511149
transform 1 0 37260 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1882_
timestamp 1644511149
transform 1 0 37260 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1883_
timestamp 1644511149
transform 1 0 36708 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1884_
timestamp 1644511149
transform 1 0 39008 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1885_
timestamp 1644511149
transform 1 0 41400 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1886_
timestamp 1644511149
transform 1 0 41216 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1887_
timestamp 1644511149
transform 1 0 42964 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1888_
timestamp 1644511149
transform 1 0 42964 0 -1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1889_
timestamp 1644511149
transform 1 0 43976 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1890_
timestamp 1644511149
transform 1 0 43240 0 -1 58752
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1891_
timestamp 1644511149
transform 1 0 44252 0 -1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1892_
timestamp 1644511149
transform 1 0 44068 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1893_
timestamp 1644511149
transform 1 0 40480 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1894_
timestamp 1644511149
transform 1 0 41124 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1895_
timestamp 1644511149
transform 1 0 35236 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1896_
timestamp 1644511149
transform 1 0 33304 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1897_
timestamp 1644511149
transform 1 0 37812 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1898_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37812 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1899_
timestamp 1644511149
transform 1 0 38916 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1900_
timestamp 1644511149
transform 1 0 28336 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _1901_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27968 0 -1 47872
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _1902_
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1903_
timestamp 1644511149
transform 1 0 38088 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1904_
timestamp 1644511149
transform 1 0 37904 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1905_
timestamp 1644511149
transform 1 0 38640 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_4  _1906_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35420 0 1 46784
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1907_
timestamp 1644511149
transform 1 0 38548 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1908_
timestamp 1644511149
transform 1 0 38272 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1909_
timestamp 1644511149
transform 1 0 38272 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1910_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27140 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1911_
timestamp 1644511149
transform 1 0 37536 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1912_
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1913_
timestamp 1644511149
transform 1 0 39008 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1914_
timestamp 1644511149
transform 1 0 38732 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1915_
timestamp 1644511149
transform 1 0 38732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1916_
timestamp 1644511149
transform 1 0 27140 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1917_
timestamp 1644511149
transform 1 0 37168 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1918_
timestamp 1644511149
transform 1 0 38088 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1919_
timestamp 1644511149
transform 1 0 38916 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1920_
timestamp 1644511149
transform 1 0 40020 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1921_
timestamp 1644511149
transform 1 0 27324 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1922_
timestamp 1644511149
transform 1 0 37352 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1923_
timestamp 1644511149
transform 1 0 38824 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1924_
timestamp 1644511149
transform 1 0 38088 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1925_
timestamp 1644511149
transform 1 0 44160 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1926_
timestamp 1644511149
transform 1 0 37904 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1927_
timestamp 1644511149
transform 1 0 37352 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1928_
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1929_
timestamp 1644511149
transform 1 0 29624 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1930_
timestamp 1644511149
transform 1 0 26404 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1931_
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1932_
timestamp 1644511149
transform 1 0 38824 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1933_
timestamp 1644511149
transform 1 0 40848 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1934_
timestamp 1644511149
transform 1 0 38916 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1935_
timestamp 1644511149
transform 1 0 39008 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1936_
timestamp 1644511149
transform 1 0 35696 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1937_
timestamp 1644511149
transform 1 0 43976 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1938_
timestamp 1644511149
transform 1 0 42872 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1939_
timestamp 1644511149
transform 1 0 27140 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1940_
timestamp 1644511149
transform 1 0 36800 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1941_
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1942_
timestamp 1644511149
transform 1 0 40664 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1943_
timestamp 1644511149
transform 1 0 40848 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1944_
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1945_
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1946_
timestamp 1644511149
transform 1 0 41492 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1947_
timestamp 1644511149
transform 1 0 42688 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1948_
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1949_
timestamp 1644511149
transform 1 0 44068 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1950_
timestamp 1644511149
transform 1 0 33488 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1951_
timestamp 1644511149
transform 1 0 36340 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1952_
timestamp 1644511149
transform 1 0 42964 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1953_
timestamp 1644511149
transform 1 0 42780 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1954_
timestamp 1644511149
transform 1 0 42780 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1955_
timestamp 1644511149
transform 1 0 33396 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1956_
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1957_
timestamp 1644511149
transform 1 0 42596 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1958_
timestamp 1644511149
transform 1 0 42504 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1959_
timestamp 1644511149
transform 1 0 45356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1960_
timestamp 1644511149
transform 1 0 45080 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1961_
timestamp 1644511149
transform 1 0 36248 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1962_
timestamp 1644511149
transform 1 0 33672 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1963_
timestamp 1644511149
transform 1 0 34592 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1964_
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1965_
timestamp 1644511149
transform 1 0 37352 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1966_
timestamp 1644511149
transform 1 0 43884 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1967_
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1968_
timestamp 1644511149
transform 1 0 42872 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1969_
timestamp 1644511149
transform 1 0 44804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1970_
timestamp 1644511149
transform 1 0 44252 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1971_
timestamp 1644511149
transform 1 0 41584 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _1972_
timestamp 1644511149
transform 1 0 33856 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1973_
timestamp 1644511149
transform 1 0 38180 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1974_
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1975_
timestamp 1644511149
transform 1 0 41308 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1976_
timestamp 1644511149
transform 1 0 45908 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1977_
timestamp 1644511149
transform 1 0 33396 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1978_
timestamp 1644511149
transform 1 0 37260 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1979_
timestamp 1644511149
transform 1 0 41032 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1980_
timestamp 1644511149
transform 1 0 41400 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1981_
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1982_
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1983_
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1984_
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1985_
timestamp 1644511149
transform 1 0 42504 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1986_
timestamp 1644511149
transform 1 0 42412 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1987_
timestamp 1644511149
transform 1 0 46092 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _1988_
timestamp 1644511149
transform 1 0 32476 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1989_
timestamp 1644511149
transform 1 0 37168 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1990_
timestamp 1644511149
transform 1 0 42504 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1991_
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1992_
timestamp 1644511149
transform 1 0 23368 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1993_
timestamp 1644511149
transform 1 0 45172 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1994_
timestamp 1644511149
transform 1 0 29256 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1995_
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1996_
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1997_
timestamp 1644511149
transform 1 0 42964 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1998_
timestamp 1644511149
transform 1 0 37628 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1999_
timestamp 1644511149
transform 1 0 41952 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2000_
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2001_
timestamp 1644511149
transform 1 0 38088 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _2002_
timestamp 1644511149
transform 1 0 27140 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _2003_
timestamp 1644511149
transform 1 0 36340 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2004_
timestamp 1644511149
transform 1 0 41032 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2005_
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2006_
timestamp 1644511149
transform 1 0 38364 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2007_
timestamp 1644511149
transform 1 0 22724 0 1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _2008_
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2009_
timestamp 1644511149
transform 1 0 22540 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _2010_
timestamp 1644511149
transform 1 0 22356 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2011_
timestamp 1644511149
transform 1 0 21528 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2012_
timestamp 1644511149
transform 1 0 20148 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _2013_
timestamp 1644511149
transform 1 0 19228 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2014_
timestamp 1644511149
transform 1 0 21160 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2015_
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _2016_
timestamp 1644511149
transform 1 0 17940 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2017_
timestamp 1644511149
transform 1 0 21804 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2018_
timestamp 1644511149
transform 1 0 23092 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2019_
timestamp 1644511149
transform 1 0 22540 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _2020_
timestamp 1644511149
transform 1 0 18400 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _2021_
timestamp 1644511149
transform 1 0 17480 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2022_
timestamp 1644511149
transform 1 0 20884 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2023_
timestamp 1644511149
transform 1 0 20608 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _2024_
timestamp 1644511149
transform 1 0 24380 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _2025_
timestamp 1644511149
transform 1 0 17848 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2026_
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2027_
timestamp 1644511149
transform 1 0 22356 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2028_
timestamp 1644511149
transform 1 0 22448 0 1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _2029_
timestamp 1644511149
transform 1 0 17572 0 -1 50048
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2030_
timestamp 1644511149
transform 1 0 22356 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _2031_
timestamp 1644511149
transform 1 0 21804 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2032_
timestamp 1644511149
transform 1 0 21712 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2033_
timestamp 1644511149
transform 1 0 20792 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _2034_
timestamp 1644511149
transform 1 0 17388 0 -1 52224
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2035_
timestamp 1644511149
transform 1 0 21528 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2036_
timestamp 1644511149
transform 1 0 22908 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _2037_
timestamp 1644511149
transform 1 0 17296 0 -1 54400
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2038_
timestamp 1644511149
transform 1 0 20792 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2039_
timestamp 1644511149
transform 1 0 24472 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2040_
timestamp 1644511149
transform 1 0 21344 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _2041_
timestamp 1644511149
transform 1 0 27968 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _2042_
timestamp 1644511149
transform 1 0 18124 0 -1 57664
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2043_
timestamp 1644511149
transform 1 0 21804 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2044_
timestamp 1644511149
transform 1 0 23644 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _2045_
timestamp 1644511149
transform 1 0 24748 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _2046_
timestamp 1644511149
transform 1 0 18584 0 -1 59840
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2047_
timestamp 1644511149
transform 1 0 21620 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2048_
timestamp 1644511149
transform 1 0 22724 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2049_
timestamp 1644511149
transform 1 0 31556 0 1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _2050_
timestamp 1644511149
transform 1 0 20792 0 1 59840
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _2051_
timestamp 1644511149
transform 1 0 32292 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2052_
timestamp 1644511149
transform 1 0 31280 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2053_
timestamp 1644511149
transform 1 0 30544 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2054_
timestamp 1644511149
transform 1 0 29532 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _2055_
timestamp 1644511149
transform 1 0 27140 0 1 59840
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2056_
timestamp 1644511149
transform 1 0 30360 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2057_
timestamp 1644511149
transform 1 0 30268 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _2058_
timestamp 1644511149
transform 1 0 27876 0 -1 58752
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2059_
timestamp 1644511149
transform 1 0 32108 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2060_
timestamp 1644511149
transform 1 0 32108 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _2061_
timestamp 1644511149
transform 1 0 28980 0 -1 56576
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2062_
timestamp 1644511149
transform 1 0 31464 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2063_
timestamp 1644511149
transform 1 0 32200 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _2064_
timestamp 1644511149
transform 1 0 28060 0 -1 53312
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2065_
timestamp 1644511149
transform 1 0 31372 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2066_
timestamp 1644511149
transform 1 0 32844 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _2067_
timestamp 1644511149
transform 1 0 29532 0 1 51136
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _2068_
timestamp 1644511149
transform 1 0 38456 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2069_
timestamp 1644511149
transform 1 0 37352 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _2070_
timestamp 1644511149
transform 1 0 40756 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2071_
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2072_
timestamp 1644511149
transform 1 0 41584 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2073_
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2074_
timestamp 1644511149
transform 1 0 39928 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2075_
timestamp 1644511149
transform 1 0 40940 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2076_
timestamp 1644511149
transform 1 0 42412 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2077_
timestamp 1644511149
transform 1 0 48392 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2078_
timestamp 1644511149
transform 1 0 46276 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2079_
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2080_
timestamp 1644511149
transform 1 0 48392 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2081_
timestamp 1644511149
transform 1 0 46736 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2082_
timestamp 1644511149
transform 1 0 48024 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2083_
timestamp 1644511149
transform 1 0 49220 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2084_
timestamp 1644511149
transform 1 0 49496 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2085_
timestamp 1644511149
transform 1 0 50876 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2086_
timestamp 1644511149
transform 1 0 50140 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2087_
timestamp 1644511149
transform 1 0 51428 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2088_
timestamp 1644511149
transform 1 0 51244 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2089_
timestamp 1644511149
transform 1 0 40020 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2090_
timestamp 1644511149
transform 1 0 45080 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2091_
timestamp 1644511149
transform 1 0 50140 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2092_
timestamp 1644511149
transform 1 0 47564 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2093_
timestamp 1644511149
transform 1 0 45724 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2094_
timestamp 1644511149
transform 1 0 50692 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2095_
timestamp 1644511149
transform 1 0 50324 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2096_
timestamp 1644511149
transform 1 0 44988 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2097_
timestamp 1644511149
transform 1 0 47564 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2098_
timestamp 1644511149
transform 1 0 48576 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2099_
timestamp 1644511149
transform 1 0 46644 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2100_
timestamp 1644511149
transform 1 0 45172 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2101_
timestamp 1644511149
transform 1 0 44160 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2102_
timestamp 1644511149
transform 1 0 40204 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2103_
timestamp 1644511149
transform 1 0 41400 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2104_
timestamp 1644511149
transform 1 0 39468 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2105_
timestamp 1644511149
transform 1 0 39008 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2106_
timestamp 1644511149
transform 1 0 30360 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2107_
timestamp 1644511149
transform 1 0 29716 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _2108_
timestamp 1644511149
transform 1 0 35512 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _2109_
timestamp 1644511149
transform 1 0 28520 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2110_
timestamp 1644511149
transform 1 0 28612 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2111_
timestamp 1644511149
transform 1 0 27416 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2112_
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2113_
timestamp 1644511149
transform 1 0 35328 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2114_
timestamp 1644511149
transform 1 0 35788 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2115_
timestamp 1644511149
transform 1 0 36156 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2116_
timestamp 1644511149
transform 1 0 35420 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2117_
timestamp 1644511149
transform 1 0 35604 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2118_
timestamp 1644511149
transform 1 0 36708 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2119_
timestamp 1644511149
transform 1 0 34776 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2120_
timestamp 1644511149
transform 1 0 31924 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2121_
timestamp 1644511149
transform 1 0 31648 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2122_
timestamp 1644511149
transform 1 0 32476 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2123_
timestamp 1644511149
transform 1 0 32384 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2124_
timestamp 1644511149
transform 1 0 29992 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2125_
timestamp 1644511149
transform 1 0 27416 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2126_
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2127_
timestamp 1644511149
transform 1 0 20976 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2128_
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2129_
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2130_
timestamp 1644511149
transform 1 0 20056 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2131_
timestamp 1644511149
transform 1 0 20240 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2132_
timestamp 1644511149
transform 1 0 19228 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2133_
timestamp 1644511149
transform 1 0 20792 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2134_
timestamp 1644511149
transform 1 0 19320 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2135_
timestamp 1644511149
transform 1 0 19412 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2136_
timestamp 1644511149
transform 1 0 19596 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2137_
timestamp 1644511149
transform 1 0 19228 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2138_
timestamp 1644511149
transform 1 0 20792 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2139_
timestamp 1644511149
transform 1 0 30360 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2140_
timestamp 1644511149
transform 1 0 29624 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2141_
timestamp 1644511149
transform 1 0 30176 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2142_
timestamp 1644511149
transform 1 0 31188 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2143_
timestamp 1644511149
transform 1 0 29900 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2144_
timestamp 1644511149
transform 1 0 30820 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2145_
timestamp 1644511149
transform 1 0 26220 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2146_
timestamp 1644511149
transform 1 0 26220 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2147_
timestamp 1644511149
transform 1 0 25852 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2148_
timestamp 1644511149
transform 1 0 25760 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2149_
timestamp 1644511149
transform 1 0 26128 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2150_
timestamp 1644511149
transform 1 0 25760 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2151_
timestamp 1644511149
transform 1 0 30176 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2152_
timestamp 1644511149
transform 1 0 30452 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2153_
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2154_
timestamp 1644511149
transform 1 0 30912 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2155_
timestamp 1644511149
transform 1 0 32384 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2156_
timestamp 1644511149
transform 1 0 32200 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2157_
timestamp 1644511149
transform 1 0 32384 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2158_
timestamp 1644511149
transform 1 0 30820 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2159_
timestamp 1644511149
transform 1 0 33212 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2160_
timestamp 1644511149
transform 1 0 33948 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2161_
timestamp 1644511149
transform 1 0 33028 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2162_
timestamp 1644511149
transform 1 0 31280 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2163_
timestamp 1644511149
transform 1 0 30912 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2164_
timestamp 1644511149
transform 1 0 22172 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _2165_
timestamp 1644511149
transform 1 0 26220 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2166_
timestamp 1644511149
transform 1 0 24104 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2167_
timestamp 1644511149
transform 1 0 18768 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2168_
timestamp 1644511149
transform 1 0 16836 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2169_
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2170_
timestamp 1644511149
transform 1 0 17388 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2171_
timestamp 1644511149
transform 1 0 16284 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2172_
timestamp 1644511149
transform 1 0 16652 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2173_
timestamp 1644511149
transform 1 0 16652 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2174_
timestamp 1644511149
transform 1 0 16560 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2175_
timestamp 1644511149
transform 1 0 15824 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2176_
timestamp 1644511149
transform 1 0 23184 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _2177_
timestamp 1644511149
transform 1 0 19688 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2178_
timestamp 1644511149
transform 1 0 21804 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2179_
timestamp 1644511149
transform 1 0 25944 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2180_
timestamp 1644511149
transform 1 0 28060 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2181_
timestamp 1644511149
transform 1 0 27508 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2182_
timestamp 1644511149
transform 1 0 29900 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2183_
timestamp 1644511149
transform 1 0 25392 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2184_
timestamp 1644511149
transform 1 0 26680 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2185_
timestamp 1644511149
transform 1 0 26128 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2186_
timestamp 1644511149
transform 1 0 26128 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2187_
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2188_
timestamp 1644511149
transform 1 0 25208 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2189_
timestamp 1644511149
transform 1 0 24748 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _2190_
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2191_
timestamp 1644511149
transform 1 0 24564 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2192_
timestamp 1644511149
transform 1 0 26128 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2193_
timestamp 1644511149
transform 1 0 29716 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2194_
timestamp 1644511149
transform 1 0 29440 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2195_
timestamp 1644511149
transform 1 0 30268 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2196_
timestamp 1644511149
transform 1 0 30452 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2197_
timestamp 1644511149
transform 1 0 30360 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2198_
timestamp 1644511149
transform 1 0 30176 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2199_
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2200_
timestamp 1644511149
transform 1 0 30912 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2201_
timestamp 1644511149
transform 1 0 23828 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2202_
timestamp 1644511149
transform 1 0 25392 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2203_
timestamp 1644511149
transform 1 0 23460 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2204_
timestamp 1644511149
transform 1 0 23920 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2205_
timestamp 1644511149
transform 1 0 23276 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2206_
timestamp 1644511149
transform 1 0 23000 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2207_
timestamp 1644511149
transform 1 0 13984 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2208_
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2209_
timestamp 1644511149
transform 1 0 12420 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2210_
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2211_
timestamp 1644511149
transform 1 0 12420 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2212_
timestamp 1644511149
transform 1 0 13984 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2213_
timestamp 1644511149
transform 1 0 29256 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2214_
timestamp 1644511149
transform 1 0 23460 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _2215_
timestamp 1644511149
transform 1 0 15548 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2216_
timestamp 1644511149
transform 1 0 15732 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2217_
timestamp 1644511149
transform 1 0 15640 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2218_
timestamp 1644511149
transform 1 0 17480 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2219_
timestamp 1644511149
transform 1 0 23552 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2220_
timestamp 1644511149
transform 1 0 24748 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2221_
timestamp 1644511149
transform 1 0 24104 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2222_
timestamp 1644511149
transform 1 0 24564 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2223_
timestamp 1644511149
transform 1 0 25024 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2224_
timestamp 1644511149
transform 1 0 23552 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2225_
timestamp 1644511149
transform 1 0 24840 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2226_
timestamp 1644511149
transform 1 0 23000 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2227_
timestamp 1644511149
transform 1 0 22264 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2228_
timestamp 1644511149
transform 1 0 22356 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2229_
timestamp 1644511149
transform 1 0 22264 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2230_
timestamp 1644511149
transform 1 0 23092 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2231_
timestamp 1644511149
transform 1 0 21896 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2232_
timestamp 1644511149
transform 1 0 30452 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2233_
timestamp 1644511149
transform 1 0 31188 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2234_
timestamp 1644511149
transform 1 0 32476 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2235_
timestamp 1644511149
transform 1 0 30912 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2236_
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2237_
timestamp 1644511149
transform 1 0 33580 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2238_
timestamp 1644511149
transform 1 0 26312 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2239_
timestamp 1644511149
transform 1 0 27048 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2240_
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2241_
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2242_
timestamp 1644511149
transform 1 0 27416 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2243_
timestamp 1644511149
transform 1 0 26128 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2244_
timestamp 1644511149
transform 1 0 32476 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2245_
timestamp 1644511149
transform 1 0 14444 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2246_
timestamp 1644511149
transform 1 0 15640 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2247_
timestamp 1644511149
transform 1 0 14720 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2248_
timestamp 1644511149
transform 1 0 14536 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2249_
timestamp 1644511149
transform 1 0 14444 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2250_
timestamp 1644511149
transform 1 0 14260 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2251_
timestamp 1644511149
transform 1 0 14168 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2252_
timestamp 1644511149
transform 1 0 14628 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2253_
timestamp 1644511149
transform 1 0 13248 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2254_
timestamp 1644511149
transform 1 0 13432 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2255_
timestamp 1644511149
transform 1 0 14168 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2256_
timestamp 1644511149
transform 1 0 13892 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2257_
timestamp 1644511149
transform 1 0 24288 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2258_
timestamp 1644511149
transform 1 0 23460 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2259_
timestamp 1644511149
transform 1 0 26220 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2260_
timestamp 1644511149
transform 1 0 26128 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2261_
timestamp 1644511149
transform 1 0 25944 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2262_
timestamp 1644511149
transform 1 0 26128 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2263_
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2264_
timestamp 1644511149
transform 1 0 36524 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _2265_
timestamp 1644511149
transform 1 0 38916 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2266_
timestamp 1644511149
transform 1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2267_
timestamp 1644511149
transform 1 0 37076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2268_
timestamp 1644511149
transform 1 0 38640 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2269_
timestamp 1644511149
transform 1 0 37628 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _2270_
timestamp 1644511149
transform 1 0 37536 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2271_
timestamp 1644511149
transform 1 0 41216 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2272_
timestamp 1644511149
transform 1 0 41216 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2273_
timestamp 1644511149
transform 1 0 43700 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2274_
timestamp 1644511149
transform 1 0 43424 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2275_
timestamp 1644511149
transform 1 0 40664 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _2276_
timestamp 1644511149
transform 1 0 43608 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2277_
timestamp 1644511149
transform 1 0 40756 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2278_
timestamp 1644511149
transform 1 0 40204 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2279_
timestamp 1644511149
transform 1 0 42136 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2280_
timestamp 1644511149
transform 1 0 43424 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2281_
timestamp 1644511149
transform 1 0 43792 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _2282_
timestamp 1644511149
transform 1 0 41584 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2283_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34868 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2284_
timestamp 1644511149
transform 1 0 36800 0 1 60928
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2285_
timestamp 1644511149
transform 1 0 33396 0 -1 62016
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2286_
timestamp 1644511149
transform 1 0 33948 0 -1 64192
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2287_
timestamp 1644511149
transform 1 0 38272 0 -1 63104
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2288_
timestamp 1644511149
transform 1 0 37904 0 1 64192
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2289_
timestamp 1644511149
transform 1 0 35144 0 1 65280
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2290_
timestamp 1644511149
transform 1 0 39836 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2291_
timestamp 1644511149
transform 1 0 42504 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2292_
timestamp 1644511149
transform 1 0 37536 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2293_
timestamp 1644511149
transform 1 0 43056 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2294_
timestamp 1644511149
transform 1 0 40112 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2295_
timestamp 1644511149
transform 1 0 32108 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2296_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32568 0 -1 47872
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2297_
timestamp 1644511149
transform 1 0 34868 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2298_
timestamp 1644511149
transform 1 0 35328 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2299_
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2300_
timestamp 1644511149
transform 1 0 37260 0 -1 48960
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2301_
timestamp 1644511149
transform 1 0 34684 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2302_
timestamp 1644511149
transform 1 0 32752 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2303_
timestamp 1644511149
transform 1 0 33580 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2304_
timestamp 1644511149
transform 1 0 33120 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2305_
timestamp 1644511149
transform 1 0 36524 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2306_
timestamp 1644511149
transform 1 0 34684 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2307_
timestamp 1644511149
transform 1 0 38088 0 -1 60928
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2308_
timestamp 1644511149
transform 1 0 39836 0 1 60928
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2309_
timestamp 1644511149
transform 1 0 37260 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2310_
timestamp 1644511149
transform 1 0 36248 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2311_
timestamp 1644511149
transform 1 0 40848 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2312_
timestamp 1644511149
transform 1 0 42872 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2313_
timestamp 1644511149
transform 1 0 44988 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2314_
timestamp 1644511149
transform 1 0 40756 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2315_
timestamp 1644511149
transform 1 0 33304 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2316_
timestamp 1644511149
transform 1 0 37904 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2317_
timestamp 1644511149
transform 1 0 39836 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2318_
timestamp 1644511149
transform 1 0 40388 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2319_
timestamp 1644511149
transform 1 0 36984 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2320_
timestamp 1644511149
transform 1 0 38824 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2321_
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2322_
timestamp 1644511149
transform 1 0 45172 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2323_
timestamp 1644511149
transform 1 0 42780 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2324_
timestamp 1644511149
transform 1 0 45448 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2325_
timestamp 1644511149
transform 1 0 45172 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2326_
timestamp 1644511149
transform 1 0 46460 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2327_
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2328_
timestamp 1644511149
transform 1 0 46736 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2329_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2330_
timestamp 1644511149
transform 1 0 46644 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2331_
timestamp 1644511149
transform 1 0 38916 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2332_
timestamp 1644511149
transform 1 0 19872 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2333_
timestamp 1644511149
transform 1 0 21068 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2334_
timestamp 1644511149
transform 1 0 22448 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2335_
timestamp 1644511149
transform 1 0 20884 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2336_
timestamp 1644511149
transform 1 0 21620 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2337_
timestamp 1644511149
transform 1 0 21804 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2338_
timestamp 1644511149
transform 1 0 23184 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2339_
timestamp 1644511149
transform 1 0 21804 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2340_
timestamp 1644511149
transform 1 0 22448 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2341_
timestamp 1644511149
transform 1 0 22448 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2342_
timestamp 1644511149
transform 1 0 31648 0 1 60928
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2343_
timestamp 1644511149
transform 1 0 29624 0 -1 62016
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2344_
timestamp 1644511149
transform 1 0 32384 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2345_
timestamp 1644511149
transform 1 0 32660 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2346_
timestamp 1644511149
transform 1 0 32108 0 -1 54400
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2347_
timestamp 1644511149
transform 1 0 37812 0 -1 52224
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2348_
timestamp 1644511149
transform 1 0 41676 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2349_
timestamp 1644511149
transform 1 0 42044 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2350_
timestamp 1644511149
transform 1 0 40020 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2351_
timestamp 1644511149
transform 1 0 39100 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2352_
timestamp 1644511149
transform 1 0 43148 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2353_
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2354_
timestamp 1644511149
transform 1 0 47564 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2355_
timestamp 1644511149
transform 1 0 48024 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2356_
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2357_
timestamp 1644511149
transform 1 0 49404 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2358_
timestamp 1644511149
transform 1 0 50140 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2359_
timestamp 1644511149
transform 1 0 51612 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2360_
timestamp 1644511149
transform 1 0 50140 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2361_
timestamp 1644511149
transform 1 0 51704 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2362_
timestamp 1644511149
transform 1 0 51520 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2363_
timestamp 1644511149
transform 1 0 49772 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2364_
timestamp 1644511149
transform 1 0 47564 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2365_
timestamp 1644511149
transform 1 0 45724 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2366_
timestamp 1644511149
transform 1 0 50508 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2367_
timestamp 1644511149
transform 1 0 50416 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2368_
timestamp 1644511149
transform 1 0 47656 0 1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2369_
timestamp 1644511149
transform 1 0 49128 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2370_
timestamp 1644511149
transform 1 0 46828 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2371_
timestamp 1644511149
transform 1 0 45172 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2372_
timestamp 1644511149
transform 1 0 43608 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2373_
timestamp 1644511149
transform 1 0 41492 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2374_
timestamp 1644511149
transform 1 0 40204 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2375_
timestamp 1644511149
transform 1 0 39468 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2376_
timestamp 1644511149
transform 1 0 30176 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2377_
timestamp 1644511149
transform 1 0 29348 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2378_
timestamp 1644511149
transform 1 0 28612 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2379_
timestamp 1644511149
transform 1 0 28704 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2380_
timestamp 1644511149
transform 1 0 26956 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2381_
timestamp 1644511149
transform 1 0 28612 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2382_
timestamp 1644511149
transform 1 0 35144 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2383_
timestamp 1644511149
transform 1 0 35512 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2384_
timestamp 1644511149
transform 1 0 35512 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2385_
timestamp 1644511149
transform 1 0 35328 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2386_
timestamp 1644511149
transform 1 0 35972 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2387_
timestamp 1644511149
transform 1 0 35512 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2388_
timestamp 1644511149
transform 1 0 34868 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2389_
timestamp 1644511149
transform 1 0 32016 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2390_
timestamp 1644511149
transform 1 0 29900 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2391_
timestamp 1644511149
transform 1 0 27600 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2392_
timestamp 1644511149
transform 1 0 25760 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2393_
timestamp 1644511149
transform 1 0 21620 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2394_
timestamp 1644511149
transform 1 0 19780 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2395_
timestamp 1644511149
transform 1 0 19872 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2396_
timestamp 1644511149
transform 1 0 20424 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2397_
timestamp 1644511149
transform 1 0 19228 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2398_
timestamp 1644511149
transform 1 0 19320 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2399_
timestamp 1644511149
transform 1 0 19596 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2400_
timestamp 1644511149
transform 1 0 19688 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2401_
timestamp 1644511149
transform 1 0 19044 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2402_
timestamp 1644511149
transform 1 0 21804 0 -1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2403_
timestamp 1644511149
transform 1 0 29348 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2404_
timestamp 1644511149
transform 1 0 30268 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2405_
timestamp 1644511149
transform 1 0 30820 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2406_
timestamp 1644511149
transform 1 0 29808 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2407_
timestamp 1644511149
transform 1 0 31096 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2408_
timestamp 1644511149
transform 1 0 27600 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2409_
timestamp 1644511149
transform 1 0 25300 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2410_
timestamp 1644511149
transform 1 0 25300 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2411_
timestamp 1644511149
transform 1 0 26220 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2412_
timestamp 1644511149
transform 1 0 25024 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2413_
timestamp 1644511149
transform 1 0 28520 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2414_
timestamp 1644511149
transform 1 0 31096 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2415_
timestamp 1644511149
transform 1 0 33120 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2416_
timestamp 1644511149
transform 1 0 32384 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2417_
timestamp 1644511149
transform 1 0 32568 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2418_
timestamp 1644511149
transform 1 0 32752 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2419_
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2420_
timestamp 1644511149
transform 1 0 32752 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2421_
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2422_
timestamp 1644511149
transform 1 0 30912 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2423_
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2424_
timestamp 1644511149
transform 1 0 24380 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2425_
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2426_
timestamp 1644511149
transform 1 0 16928 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2427_
timestamp 1644511149
transform 1 0 16468 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2428_
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2429_
timestamp 1644511149
transform 1 0 16284 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2430_
timestamp 1644511149
transform 1 0 16744 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2431_
timestamp 1644511149
transform 1 0 16928 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2432_
timestamp 1644511149
transform 1 0 16652 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2433_
timestamp 1644511149
transform 1 0 19228 0 -1 62016
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2434_
timestamp 1644511149
transform 1 0 21160 0 1 60928
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2435_
timestamp 1644511149
transform 1 0 26220 0 1 62016
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2436_
timestamp 1644511149
transform 1 0 27508 0 -1 62016
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2437_
timestamp 1644511149
transform 1 0 27140 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2438_
timestamp 1644511149
transform 1 0 26772 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2439_
timestamp 1644511149
transform 1 0 26956 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2440_
timestamp 1644511149
transform 1 0 26404 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2441_
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2442_
timestamp 1644511149
transform 1 0 24196 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2443_
timestamp 1644511149
transform 1 0 24380 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2444_
timestamp 1644511149
transform 1 0 24656 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2445_
timestamp 1644511149
transform 1 0 25024 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2446_
timestamp 1644511149
transform 1 0 30176 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2447_
timestamp 1644511149
transform 1 0 29716 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2448_
timestamp 1644511149
transform 1 0 30544 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2449_
timestamp 1644511149
transform 1 0 30176 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2450_
timestamp 1644511149
transform 1 0 30912 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2451_
timestamp 1644511149
transform 1 0 31372 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2452_
timestamp 1644511149
transform 1 0 31280 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2453_
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2454_
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2455_
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2456_
timestamp 1644511149
transform 1 0 23276 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2457_
timestamp 1644511149
transform 1 0 16744 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2458_
timestamp 1644511149
transform 1 0 12696 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2459_
timestamp 1644511149
transform 1 0 12512 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2460_
timestamp 1644511149
transform 1 0 12144 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2461_
timestamp 1644511149
transform 1 0 12420 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2462_
timestamp 1644511149
transform 1 0 14352 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2463_
timestamp 1644511149
transform 1 0 15548 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2464_
timestamp 1644511149
transform 1 0 16468 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2465_
timestamp 1644511149
transform 1 0 15548 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2466_
timestamp 1644511149
transform 1 0 17388 0 -1 60928
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2467_
timestamp 1644511149
transform 1 0 24380 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2468_
timestamp 1644511149
transform 1 0 24840 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2469_
timestamp 1644511149
transform 1 0 24472 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2470_
timestamp 1644511149
transform 1 0 24840 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2471_
timestamp 1644511149
transform 1 0 24840 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2472_
timestamp 1644511149
transform 1 0 25484 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2473_
timestamp 1644511149
transform 1 0 22264 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2474_
timestamp 1644511149
transform 1 0 22448 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2475_
timestamp 1644511149
transform 1 0 22356 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2476_
timestamp 1644511149
transform 1 0 23460 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2477_
timestamp 1644511149
transform 1 0 21804 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2478_
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2479_
timestamp 1644511149
transform 1 0 32660 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2480_
timestamp 1644511149
transform 1 0 31096 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2481_
timestamp 1644511149
transform 1 0 34592 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2482_
timestamp 1644511149
transform 1 0 33672 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2483_
timestamp 1644511149
transform 1 0 27048 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2484_
timestamp 1644511149
transform 1 0 29256 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2485_
timestamp 1644511149
transform 1 0 29900 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2486_
timestamp 1644511149
transform 1 0 27600 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2487_
timestamp 1644511149
transform 1 0 26220 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2488_
timestamp 1644511149
transform 1 0 22264 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2489_
timestamp 1644511149
transform 1 0 14720 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2490_
timestamp 1644511149
transform 1 0 14628 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2491_
timestamp 1644511149
transform 1 0 14536 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2492_
timestamp 1644511149
transform 1 0 14168 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2493_
timestamp 1644511149
transform 1 0 14260 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2494_
timestamp 1644511149
transform 1 0 13524 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2495_
timestamp 1644511149
transform 1 0 14168 0 -1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2496_
timestamp 1644511149
transform 1 0 14352 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2497_
timestamp 1644511149
transform 1 0 14076 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2498_
timestamp 1644511149
transform 1 0 22816 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2499_
timestamp 1644511149
transform 1 0 26956 0 -1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2500_
timestamp 1644511149
transform 1 0 26680 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2501_
timestamp 1644511149
transform 1 0 26128 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2502_
timestamp 1644511149
transform 1 0 26956 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2503_
timestamp 1644511149
transform 1 0 30176 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2504_
timestamp 1644511149
transform 1 0 38824 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2505_
timestamp 1644511149
transform 1 0 37904 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2506_
timestamp 1644511149
transform 1 0 37812 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2507_
timestamp 1644511149
transform 1 0 39284 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2508_
timestamp 1644511149
transform 1 0 37536 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2509_
timestamp 1644511149
transform 1 0 40480 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2510_
timestamp 1644511149
transform 1 0 41308 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2511_
timestamp 1644511149
transform 1 0 44068 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2512_
timestamp 1644511149
transform 1 0 43608 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2513_
timestamp 1644511149
transform 1 0 43424 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2514_
timestamp 1644511149
transform 1 0 40480 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2515_
timestamp 1644511149
transform 1 0 39928 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2516_
timestamp 1644511149
transform 1 0 42872 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2517_
timestamp 1644511149
transform 1 0 43792 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2518_
timestamp 1644511149
transform 1 0 43792 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2519_
timestamp 1644511149
transform 1 0 41124 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _2520__38 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2521__39
timestamp 1644511149
transform 1 0 4416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2522__40
timestamp 1644511149
transform 1 0 67436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2523__41
timestamp 1644511149
transform 1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2524__42
timestamp 1644511149
transform 1 0 1472 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2525__43
timestamp 1644511149
transform 1 0 36432 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2526__44
timestamp 1644511149
transform 1 0 67436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2527__45
timestamp 1644511149
transform 1 0 67712 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2528__46
timestamp 1644511149
transform 1 0 2300 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2529__47
timestamp 1644511149
transform 1 0 67896 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2530__48
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2531__49
timestamp 1644511149
transform 1 0 38180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2532__50
timestamp 1644511149
transform 1 0 1656 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2533__51
timestamp 1644511149
transform 1 0 42688 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2534__52
timestamp 1644511149
transform 1 0 64860 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2535__53
timestamp 1644511149
transform 1 0 1748 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2536__54
timestamp 1644511149
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2537__55
timestamp 1644511149
transform 1 0 24656 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2538__56
timestamp 1644511149
transform 1 0 67712 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2539__57
timestamp 1644511149
transform 1 0 60444 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2540__58
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2541__59
timestamp 1644511149
transform 1 0 60720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2542__60
timestamp 1644511149
transform 1 0 64216 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2543__61
timestamp 1644511149
transform 1 0 45908 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2544__62
timestamp 1644511149
transform 1 0 67436 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2545__63
timestamp 1644511149
transform 1 0 1748 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2546__64
timestamp 1644511149
transform 1 0 66792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2547__65
timestamp 1644511149
transform 1 0 67712 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2548__66
timestamp 1644511149
transform 1 0 41216 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2549__67
timestamp 1644511149
transform 1 0 50508 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2550__68
timestamp 1644511149
transform 1 0 1472 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2551__69
timestamp 1644511149
transform 1 0 45264 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2552__70
timestamp 1644511149
transform 1 0 16652 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2553__71
timestamp 1644511149
transform 1 0 27140 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2554__72
timestamp 1644511149
transform 1 0 37352 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2555__73
timestamp 1644511149
transform 1 0 66700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2556__74
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2557__75
timestamp 1644511149
transform 1 0 67712 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2558__76
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2559__77
timestamp 1644511149
transform 1 0 66240 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2560__78
timestamp 1644511149
transform 1 0 1564 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2561__79
timestamp 1644511149
transform 1 0 11500 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2562__80
timestamp 1644511149
transform 1 0 67712 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2563__81
timestamp 1644511149
transform 1 0 1656 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2564__82
timestamp 1644511149
transform 1 0 6348 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2565__83
timestamp 1644511149
transform 1 0 66792 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2566__84
timestamp 1644511149
transform 1 0 67712 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2567__85
timestamp 1644511149
transform 1 0 1840 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2568__86
timestamp 1644511149
transform 1 0 48760 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2569__87
timestamp 1644511149
transform 1 0 61916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2570__88
timestamp 1644511149
transform 1 0 52716 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2571__89
timestamp 1644511149
transform 1 0 67712 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2572__90
timestamp 1644511149
transform 1 0 67436 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2573__91
timestamp 1644511149
transform 1 0 67068 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2574__92
timestamp 1644511149
transform 1 0 3220 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2575__93
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2576__94
timestamp 1644511149
transform 1 0 62008 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2577__95
timestamp 1644511149
transform 1 0 1564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2578__96
timestamp 1644511149
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2579__97
timestamp 1644511149
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2580__98
timestamp 1644511149
transform 1 0 66792 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2581__99
timestamp 1644511149
transform 1 0 56304 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2582__100
timestamp 1644511149
transform 1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2583__101
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2584__102
timestamp 1644511149
transform 1 0 66792 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2585__103
timestamp 1644511149
transform 1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2586__104
timestamp 1644511149
transform 1 0 1840 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2587__105
timestamp 1644511149
transform 1 0 31004 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2588__106
timestamp 1644511149
transform 1 0 4600 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2589__107
timestamp 1644511149
transform 1 0 64860 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2590__108
timestamp 1644511149
transform 1 0 38824 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2591__109
timestamp 1644511149
transform 1 0 67712 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2592__110
timestamp 1644511149
transform 1 0 67436 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2593__111
timestamp 1644511149
transform 1 0 1932 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2594__112
timestamp 1644511149
transform 1 0 57132 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2595__113
timestamp 1644511149
transform 1 0 67712 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2596_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32292 0 1 55488
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2597_
timestamp 1644511149
transform 1 0 37168 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2598_
timestamp 1644511149
transform 1 0 49864 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2599_
timestamp 1644511149
transform 1 0 41308 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2600_
timestamp 1644511149
transform 1 0 23000 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2601_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2602_
timestamp 1644511149
transform 1 0 40020 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2603_
timestamp 1644511149
transform 1 0 46736 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2604_
timestamp 1644511149
transform 1 0 44068 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2605_
timestamp 1644511149
transform 1 0 47472 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2606_
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2607_
timestamp 1644511149
transform 1 0 47932 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2608_
timestamp 1644511149
transform 1 0 45816 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2609_
timestamp 1644511149
transform 1 0 48760 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2610_
timestamp 1644511149
transform 1 0 48576 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2611_
timestamp 1644511149
transform 1 0 48760 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2612_
timestamp 1644511149
transform 1 0 48668 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2613_
timestamp 1644511149
transform 1 0 19320 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2614_
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2615_
timestamp 1644511149
transform 1 0 23828 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2616_
timestamp 1644511149
transform 1 0 19412 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2617_
timestamp 1644511149
transform 1 0 22448 0 -1 50048
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2618_
timestamp 1644511149
transform 1 0 22724 0 -1 62016
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2619_
timestamp 1644511149
transform 1 0 29072 0 -1 63104
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2620_
timestamp 1644511149
transform 1 0 21988 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2621_
timestamp 1644511149
transform 1 0 24380 0 1 50048
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2622_
timestamp 1644511149
transform 1 0 24380 0 1 57664
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2623_
timestamp 1644511149
transform 1 0 32936 0 -1 63104
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2624_
timestamp 1644511149
transform 1 0 30360 0 1 62016
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2625_
timestamp 1644511149
transform 1 0 33672 0 -1 57664
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2626_
timestamp 1644511149
transform 1 0 33764 0 -1 59840
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2627_
timestamp 1644511149
transform 1 0 6348 0 -1 54400
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2628_
timestamp 1644511149
transform 1 0 66240 0 1 51136
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2629_
timestamp 1644511149
transform 1 0 1380 0 1 66368
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2630_
timestamp 1644511149
transform 1 0 4416 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2631_
timestamp 1644511149
transform 1 0 66240 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2632_
timestamp 1644511149
transform 1 0 10396 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2633_
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2634_
timestamp 1644511149
transform 1 0 36248 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2635_
timestamp 1644511149
transform 1 0 66240 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2636_
timestamp 1644511149
transform 1 0 65780 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2637_
timestamp 1644511149
transform 1 0 1380 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2638_
timestamp 1644511149
transform 1 0 65780 0 -1 60928
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2639_
timestamp 1644511149
transform 1 0 1564 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2640_
timestamp 1644511149
transform 1 0 38088 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2641_
timestamp 1644511149
transform 1 0 1656 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2642_
timestamp 1644511149
transform 1 0 42596 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2643_
timestamp 1644511149
transform 1 0 66240 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2644_
timestamp 1644511149
transform 1 0 1656 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2645_
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2646_
timestamp 1644511149
transform 1 0 24656 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2647_
timestamp 1644511149
transform 1 0 65780 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2648_
timestamp 1644511149
transform 1 0 60444 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2649_
timestamp 1644511149
transform 1 0 1656 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2650_
timestamp 1644511149
transform 1 0 60628 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2651_
timestamp 1644511149
transform 1 0 65504 0 -1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2652_
timestamp 1644511149
transform 1 0 46368 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2653_
timestamp 1644511149
transform 1 0 66240 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2654_
timestamp 1644511149
transform 1 0 1380 0 1 53312
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2655_
timestamp 1644511149
transform 1 0 65780 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2656_
timestamp 1644511149
transform 1 0 65780 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2657_
timestamp 1644511149
transform 1 0 40296 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2658_
timestamp 1644511149
transform 1 0 50416 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2659_
timestamp 1644511149
transform 1 0 1748 0 -1 65280
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2660_
timestamp 1644511149
transform 1 0 45172 0 -1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2661_
timestamp 1644511149
transform 1 0 16100 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2662_
timestamp 1644511149
transform 1 0 27048 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2663_
timestamp 1644511149
transform 1 0 37260 0 -1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2664_
timestamp 1644511149
transform 1 0 65780 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2665_
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2666_
timestamp 1644511149
transform 1 0 65780 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2667_
timestamp 1644511149
transform 1 0 46184 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2668_
timestamp 1644511149
transform 1 0 65780 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2669_
timestamp 1644511149
transform 1 0 1380 0 1 52224
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2670_
timestamp 1644511149
transform 1 0 11040 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2671_
timestamp 1644511149
transform 1 0 65780 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2672_
timestamp 1644511149
transform 1 0 1656 0 -1 59840
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2673_
timestamp 1644511149
transform 1 0 5980 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2674_
timestamp 1644511149
transform 1 0 65780 0 -1 67456
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2675_
timestamp 1644511149
transform 1 0 65780 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2676_
timestamp 1644511149
transform 1 0 1840 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2677_
timestamp 1644511149
transform 1 0 49588 0 -1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2678_
timestamp 1644511149
transform 1 0 61916 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2679_
timestamp 1644511149
transform 1 0 52716 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2680_
timestamp 1644511149
transform 1 0 66240 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2681_
timestamp 1644511149
transform 1 0 66240 0 1 57664
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2682_
timestamp 1644511149
transform 1 0 65780 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2683_
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2684_
timestamp 1644511149
transform 1 0 34040 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2685_
timestamp 1644511149
transform 1 0 62744 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2686_
timestamp 1644511149
transform 1 0 1564 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2687_
timestamp 1644511149
transform 1 0 3864 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2688_
timestamp 1644511149
transform 1 0 19320 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2689_
timestamp 1644511149
transform 1 0 65780 0 -1 66368
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2690_
timestamp 1644511149
transform 1 0 56212 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2691_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2692_
timestamp 1644511149
transform 1 0 21896 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2693_
timestamp 1644511149
transform 1 0 66240 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2694_
timestamp 1644511149
transform 1 0 44620 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2695_
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2696_
timestamp 1644511149
transform 1 0 31004 0 1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2697_
timestamp 1644511149
transform 1 0 4508 0 1 67456
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2698_
timestamp 1644511149
transform 1 0 65780 0 -1 69632
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2699_
timestamp 1644511149
transform 1 0 39560 0 -1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2700_
timestamp 1644511149
transform 1 0 65780 0 -1 62016
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2701_
timestamp 1644511149
transform 1 0 66240 0 1 63104
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2702_
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2703_
timestamp 1644511149
transform 1 0 57868 0 -1 68544
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2704_
timestamp 1644511149
transform 1 0 65780 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34040 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 38088 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 35052 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 34684 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 40296 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 29624 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 37996 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 32016 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 34592 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 41400 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 28704 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 30728 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 39468 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 38640 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1644511149
transform 1 0 1380 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 67620 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 1644511149
transform 1 0 67620 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1644511149
transform 1 0 67160 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1644511149
transform 1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1644511149
transform 1 0 27140 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1644511149
transform 1 0 67804 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1644511149
transform 1 0 35512 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 32292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1644511149
transform 1 0 67804 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input12
timestamp 1644511149
transform 1 0 67160 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 1644511149
transform 1 0 1380 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 1644511149
transform 1 0 67160 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1644511149
transform 1 0 1380 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1644511149
transform 1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input18
timestamp 1644511149
transform 1 0 65596 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1644511149
transform 1 0 20700 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1644511149
transform 1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1644511149
transform 1 0 19596 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1644511149
transform 1 0 7820 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input27
timestamp 1644511149
transform 1 0 67620 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input28
timestamp 1644511149
transform 1 0 42780 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input29
timestamp 1644511149
transform 1 0 67620 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input31
timestamp 1644511149
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1644511149
transform 1 0 14444 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input33
timestamp 1644511149
transform 1 0 56120 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1644511149
transform 1 0 1748 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1644511149
transform 1 0 55476 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input36
timestamp 1644511149
transform 1 0 1748 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input37
timestamp 1644511149
transform 1 0 67160 0 -1 34816
box -38 -48 590 592
<< labels >>
rlabel metal3 s 0 71348 800 71588 6 active
port 0 nsew signal input
rlabel metal3 s 69200 22388 70000 22628 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 52154 0 52266 800 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 54730 0 54842 800 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 69200 11508 70000 11748 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 69200 8788 70000 9028 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 0 10148 800 10388 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 69200 36668 70000 36908 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 69200 27148 70000 27388 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 57306 0 57418 800 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 71200 21998 72000 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 69200 1988 70000 2228 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 69200 52308 70000 52548 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 9006 71200 9118 72000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 59238 71200 59350 72000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 64390 71200 64502 72000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 32834 71200 32946 72000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 53442 0 53554 800 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 12870 71200 12982 72000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 1278 71200 1390 72000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 18022 71200 18134 72000 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 69200 3348 70000 3588 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 69200 24428 70000 24668 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 64548 800 64788 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 69200 48228 70000 48468 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 59882 0 59994 800 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 0 57748 800 57988 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 30902 0 31014 800 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 58594 0 58706 800 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 0 14228 800 14468 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 io_oeb[0]
port 39 nsew signal bidirectional
rlabel metal2 s 50222 71200 50334 72000 6 io_oeb[10]
port 40 nsew signal bidirectional
rlabel metal2 s 62458 0 62570 800 6 io_oeb[11]
port 41 nsew signal bidirectional
rlabel metal2 s 52798 71200 52910 72000 6 io_oeb[12]
port 42 nsew signal bidirectional
rlabel metal3 s 69200 43468 70000 43708 6 io_oeb[13]
port 43 nsew signal bidirectional
rlabel metal3 s 69200 57748 70000 57988 6 io_oeb[14]
port 44 nsew signal bidirectional
rlabel metal3 s 69200 42108 70000 42348 6 io_oeb[15]
port 45 nsew signal bidirectional
rlabel metal3 s 0 23748 800 23988 6 io_oeb[16]
port 46 nsew signal bidirectional
rlabel metal2 s 34766 0 34878 800 6 io_oeb[17]
port 47 nsew signal bidirectional
rlabel metal2 s 63102 71200 63214 72000 6 io_oeb[18]
port 48 nsew signal bidirectional
rlabel metal3 s 0 12868 800 13108 6 io_oeb[19]
port 49 nsew signal bidirectional
rlabel metal3 s 69200 4708 70000 4948 6 io_oeb[1]
port 50 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 io_oeb[20]
port 51 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 io_oeb[21]
port 52 nsew signal bidirectional
rlabel metal3 s 69200 65908 70000 66148 6 io_oeb[22]
port 53 nsew signal bidirectional
rlabel metal2 s 56662 71200 56774 72000 6 io_oeb[23]
port 54 nsew signal bidirectional
rlabel metal2 s 5786 0 5898 800 6 io_oeb[24]
port 55 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 io_oeb[25]
port 56 nsew signal bidirectional
rlabel metal3 s 69200 40748 70000 40988 6 io_oeb[26]
port 57 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 io_oeb[27]
port 58 nsew signal bidirectional
rlabel metal3 s 0 22388 800 22628 6 io_oeb[28]
port 59 nsew signal bidirectional
rlabel metal2 s 31546 71200 31658 72000 6 io_oeb[29]
port 60 nsew signal bidirectional
rlabel metal3 s 0 52308 800 52548 6 io_oeb[2]
port 61 nsew signal bidirectional
rlabel metal2 s 5142 71200 5254 72000 6 io_oeb[30]
port 62 nsew signal bidirectional
rlabel metal2 s 68254 71200 68366 72000 6 io_oeb[31]
port 63 nsew signal bidirectional
rlabel metal2 s 39274 71200 39386 72000 6 io_oeb[32]
port 64 nsew signal bidirectional
rlabel metal3 s 69200 61828 70000 62068 6 io_oeb[33]
port 65 nsew signal bidirectional
rlabel metal3 s 69200 63188 70000 63428 6 io_oeb[34]
port 66 nsew signal bidirectional
rlabel metal3 s 0 35308 800 35548 6 io_oeb[35]
port 67 nsew signal bidirectional
rlabel metal2 s 57950 71200 58062 72000 6 io_oeb[36]
port 68 nsew signal bidirectional
rlabel metal3 s 69200 46188 70000 46428 6 io_oeb[37]
port 69 nsew signal bidirectional
rlabel metal2 s 11582 71200 11694 72000 6 io_oeb[3]
port 70 nsew signal bidirectional
rlabel metal3 s 69200 21028 70000 21268 6 io_oeb[4]
port 71 nsew signal bidirectional
rlabel metal3 s 0 59108 800 59348 6 io_oeb[5]
port 72 nsew signal bidirectional
rlabel metal2 s 6430 71200 6542 72000 6 io_oeb[6]
port 73 nsew signal bidirectional
rlabel metal3 s 69200 67268 70000 67508 6 io_oeb[7]
port 74 nsew signal bidirectional
rlabel metal3 s 69200 35308 70000 35548 6 io_oeb[8]
port 75 nsew signal bidirectional
rlabel metal3 s 0 29868 800 30108 6 io_oeb[9]
port 76 nsew signal bidirectional
rlabel metal3 s 0 67268 800 67508 6 io_out[0]
port 77 nsew signal bidirectional
rlabel metal3 s 0 1988 800 2228 6 io_out[10]
port 78 nsew signal bidirectional
rlabel metal2 s 38630 0 38742 800 6 io_out[11]
port 79 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 io_out[12]
port 80 nsew signal bidirectional
rlabel metal2 s 43138 71200 43250 72000 6 io_out[13]
port 81 nsew signal bidirectional
rlabel metal2 s 69542 71200 69654 72000 6 io_out[14]
port 82 nsew signal bidirectional
rlabel metal3 s 0 47548 800 47788 6 io_out[15]
port 83 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 io_out[16]
port 84 nsew signal bidirectional
rlabel metal2 s 25106 71200 25218 72000 6 io_out[17]
port 85 nsew signal bidirectional
rlabel metal3 s 69200 16948 70000 17188 6 io_out[18]
port 86 nsew signal bidirectional
rlabel metal2 s 60526 71200 60638 72000 6 io_out[19]
port 87 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 io_out[1]
port 88 nsew signal bidirectional
rlabel metal3 s 0 25788 800 26028 6 io_out[20]
port 89 nsew signal bidirectional
rlabel metal2 s 61170 0 61282 800 6 io_out[21]
port 90 nsew signal bidirectional
rlabel metal2 s 66966 71200 67078 72000 6 io_out[22]
port 91 nsew signal bidirectional
rlabel metal2 s 47002 71200 47114 72000 6 io_out[23]
port 92 nsew signal bidirectional
rlabel metal3 s 69200 44828 70000 45068 6 io_out[24]
port 93 nsew signal bidirectional
rlabel metal3 s 0 53668 800 53908 6 io_out[25]
port 94 nsew signal bidirectional
rlabel metal2 s 69542 0 69654 800 6 io_out[26]
port 95 nsew signal bidirectional
rlabel metal3 s 69200 31228 70000 31468 6 io_out[27]
port 96 nsew signal bidirectional
rlabel metal2 s 41850 71200 41962 72000 6 io_out[28]
port 97 nsew signal bidirectional
rlabel metal2 s 51510 71200 51622 72000 6 io_out[29]
port 98 nsew signal bidirectional
rlabel metal3 s 69200 23068 70000 23308 6 io_out[2]
port 99 nsew signal bidirectional
rlabel metal3 s 0 4708 800 4948 6 io_out[30]
port 100 nsew signal bidirectional
rlabel metal2 s 45714 71200 45826 72000 6 io_out[31]
port 101 nsew signal bidirectional
rlabel metal2 s 16734 71200 16846 72000 6 io_out[32]
port 102 nsew signal bidirectional
rlabel metal2 s 27682 71200 27794 72000 6 io_out[33]
port 103 nsew signal bidirectional
rlabel metal2 s 37986 71200 38098 72000 6 io_out[34]
port 104 nsew signal bidirectional
rlabel metal2 s 68898 0 69010 800 6 io_out[35]
port 105 nsew signal bidirectional
rlabel metal3 s 0 15588 800 15828 6 io_out[36]
port 106 nsew signal bidirectional
rlabel metal3 s 69200 6068 70000 6308 6 io_out[37]
port 107 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 io_out[3]
port 108 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 io_out[4]
port 109 nsew signal bidirectional
rlabel metal2 s 36698 71200 36810 72000 6 io_out[5]
port 110 nsew signal bidirectional
rlabel metal3 s 69200 32588 70000 32828 6 io_out[6]
port 111 nsew signal bidirectional
rlabel metal3 s 69200 14228 70000 14468 6 io_out[7]
port 112 nsew signal bidirectional
rlabel metal3 s 0 68628 800 68868 6 io_out[8]
port 113 nsew signal bidirectional
rlabel metal3 s 69200 60468 70000 60708 6 io_out[9]
port 114 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 69680 6 vccd1
port 115 nsew power input
rlabel metal4 s 34928 2128 35248 69680 6 vccd1
port 115 nsew power input
rlabel metal4 s 65648 2128 65968 69680 6 vccd1
port 115 nsew power input
rlabel metal4 s 19568 2128 19888 69680 6 vssd1
port 116 nsew ground input
rlabel metal4 s 50288 2128 50608 69680 6 vssd1
port 116 nsew ground input
rlabel metal2 s 23174 71200 23286 72000 6 wb_clk_i
port 117 nsew signal input
rlabel metal3 s 69200 69988 70000 70228 6 wb_rst_i
port 118 nsew signal input
rlabel metal3 s 0 50948 800 51188 6 wbs_ack_o
port 119 nsew signal bidirectional
rlabel metal3 s 69200 47548 70000 47788 6 wbs_adr_i[0]
port 120 nsew signal input
rlabel metal3 s 69200 59108 70000 59348 6 wbs_adr_i[10]
port 121 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 wbs_adr_i[11]
port 122 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 wbs_adr_i[12]
port 123 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 wbs_adr_i[13]
port 124 nsew signal input
rlabel metal3 s 69200 18308 70000 18548 6 wbs_adr_i[14]
port 125 nsew signal input
rlabel metal2 s 35410 71200 35522 72000 6 wbs_adr_i[15]
port 126 nsew signal input
rlabel metal2 s 32190 0 32302 800 6 wbs_adr_i[16]
port 127 nsew signal input
rlabel metal3 s 69200 12868 70000 13108 6 wbs_adr_i[17]
port 128 nsew signal input
rlabel metal2 s 67610 0 67722 800 6 wbs_adr_i[18]
port 129 nsew signal input
rlabel metal3 s 0 63188 800 63428 6 wbs_adr_i[19]
port 130 nsew signal input
rlabel metal3 s 0 46188 800 46428 6 wbs_adr_i[1]
port 131 nsew signal input
rlabel metal3 s 69200 39388 70000 39628 6 wbs_adr_i[20]
port 132 nsew signal input
rlabel metal3 s 0 56388 800 56628 6 wbs_adr_i[21]
port 133 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 wbs_adr_i[22]
port 134 nsew signal input
rlabel metal2 s 65034 0 65146 800 6 wbs_adr_i[23]
port 135 nsew signal input
rlabel metal2 s 20598 71200 20710 72000 6 wbs_adr_i[24]
port 136 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 wbs_adr_i[25]
port 137 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 wbs_adr_i[26]
port 138 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 wbs_adr_i[27]
port 139 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 wbs_adr_i[28]
port 140 nsew signal input
rlabel metal2 s 19310 71200 19422 72000 6 wbs_adr_i[29]
port 141 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 wbs_adr_i[2]
port 142 nsew signal input
rlabel metal2 s 7718 71200 7830 72000 6 wbs_adr_i[30]
port 143 nsew signal input
rlabel metal3 s 69200 7428 70000 7668 6 wbs_adr_i[31]
port 144 nsew signal input
rlabel metal2 s 42494 0 42606 800 6 wbs_adr_i[3]
port 145 nsew signal input
rlabel metal3 s 69200 56388 70000 56628 6 wbs_adr_i[4]
port 146 nsew signal input
rlabel metal3 s 0 7428 800 7668 6 wbs_adr_i[5]
port 147 nsew signal input
rlabel metal2 s 17378 0 17490 800 6 wbs_adr_i[6]
port 148 nsew signal input
rlabel metal2 s 14158 71200 14270 72000 6 wbs_adr_i[7]
port 149 nsew signal input
rlabel metal2 s 56018 0 56130 800 6 wbs_adr_i[8]
port 150 nsew signal input
rlabel metal3 s 0 43468 800 43708 6 wbs_adr_i[9]
port 151 nsew signal input
rlabel metal2 s 55374 71200 55486 72000 6 wbs_cyc_i
port 152 nsew signal input
rlabel metal2 s 634 71200 746 72000 6 wbs_dat_i[0]
port 153 nsew signal input
rlabel metal2 s 15446 71200 15558 72000 6 wbs_dat_i[10]
port 154 nsew signal input
rlabel metal2 s 26394 71200 26506 72000 6 wbs_dat_i[11]
port 155 nsew signal input
rlabel metal2 s 23818 71200 23930 72000 6 wbs_dat_i[12]
port 156 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 wbs_dat_i[13]
port 157 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 wbs_dat_i[14]
port 158 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 wbs_dat_i[15]
port 159 nsew signal input
rlabel metal2 s 33478 0 33590 800 6 wbs_dat_i[16]
port 160 nsew signal input
rlabel metal3 s 69200 68628 70000 68868 6 wbs_dat_i[17]
port 161 nsew signal input
rlabel metal2 s 2566 71200 2678 72000 6 wbs_dat_i[18]
port 162 nsew signal input
rlabel metal2 s 34122 71200 34234 72000 6 wbs_dat_i[19]
port 163 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 wbs_dat_i[1]
port 164 nsew signal input
rlabel metal3 s 69200 25788 70000 26028 6 wbs_dat_i[20]
port 165 nsew signal input
rlabel metal3 s 69200 53668 70000 53908 6 wbs_dat_i[21]
port 166 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 wbs_dat_i[22]
port 167 nsew signal input
rlabel metal3 s 69200 38028 70000 38268 6 wbs_dat_i[23]
port 168 nsew signal input
rlabel metal3 s 0 61828 800 62068 6 wbs_dat_i[24]
port 169 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 wbs_dat_i[25]
port 170 nsew signal input
rlabel metal3 s 69200 64548 70000 64788 6 wbs_dat_i[26]
port 171 nsew signal input
rlabel metal2 s 40562 71200 40674 72000 6 wbs_dat_i[27]
port 172 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 wbs_dat_i[28]
port 173 nsew signal input
rlabel metal3 s 69200 28508 70000 28748 6 wbs_dat_i[29]
port 174 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 wbs_dat_i[2]
port 175 nsew signal input
rlabel metal3 s 69200 10148 70000 10388 6 wbs_dat_i[30]
port 176 nsew signal input
rlabel metal3 s 0 65908 800 66148 6 wbs_dat_i[31]
port 177 nsew signal input
rlabel metal2 s 63746 0 63858 800 6 wbs_dat_i[3]
port 178 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 wbs_dat_i[4]
port 179 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 wbs_dat_i[5]
port 180 nsew signal input
rlabel metal3 s 69200 19668 70000 19908 6 wbs_dat_i[6]
port 181 nsew signal input
rlabel metal3 s 69200 71348 70000 71588 6 wbs_dat_i[7]
port 182 nsew signal input
rlabel metal3 s 0 18308 800 18548 6 wbs_dat_i[8]
port 183 nsew signal input
rlabel metal2 s 66322 0 66434 800 6 wbs_dat_i[9]
port 184 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 wbs_dat_o[0]
port 185 nsew signal bidirectional
rlabel metal3 s 69200 29868 70000 30108 6 wbs_dat_o[10]
port 186 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 wbs_dat_o[11]
port 187 nsew signal bidirectional
rlabel metal3 s 69200 55028 70000 55268 6 wbs_dat_o[12]
port 188 nsew signal bidirectional
rlabel metal2 s 65678 71200 65790 72000 6 wbs_dat_o[13]
port 189 nsew signal bidirectional
rlabel metal3 s 69200 628 70000 868 6 wbs_dat_o[14]
port 190 nsew signal bidirectional
rlabel metal2 s 61814 71200 61926 72000 6 wbs_dat_o[15]
port 191 nsew signal bidirectional
rlabel metal3 s 0 38028 800 38268 6 wbs_dat_o[16]
port 192 nsew signal bidirectional
rlabel metal3 s 0 40748 800 40988 6 wbs_dat_o[17]
port 193 nsew signal bidirectional
rlabel metal2 s 43782 0 43894 800 6 wbs_dat_o[18]
port 194 nsew signal bidirectional
rlabel metal2 s -10 0 102 800 6 wbs_dat_o[19]
port 195 nsew signal bidirectional
rlabel metal2 s 50866 0 50978 800 6 wbs_dat_o[1]
port 196 nsew signal bidirectional
rlabel metal3 s 0 49588 800 49828 6 wbs_dat_o[20]
port 197 nsew signal bidirectional
rlabel metal2 s 3854 71200 3966 72000 6 wbs_dat_o[21]
port 198 nsew signal bidirectional
rlabel metal2 s 30258 71200 30370 72000 6 wbs_dat_o[22]
port 199 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 wbs_dat_o[23]
port 200 nsew signal bidirectional
rlabel metal2 s 13514 0 13626 800 6 wbs_dat_o[24]
port 201 nsew signal bidirectional
rlabel metal2 s 4498 0 4610 800 6 wbs_dat_o[25]
port 202 nsew signal bidirectional
rlabel metal2 s 44426 71200 44538 72000 6 wbs_dat_o[26]
port 203 nsew signal bidirectional
rlabel metal2 s 28970 71200 29082 72000 6 wbs_dat_o[27]
port 204 nsew signal bidirectional
rlabel metal2 s 36054 0 36166 800 6 wbs_dat_o[28]
port 205 nsew signal bidirectional
rlabel metal2 s 54086 71200 54198 72000 6 wbs_dat_o[29]
port 206 nsew signal bidirectional
rlabel metal3 s 69200 15588 70000 15828 6 wbs_dat_o[2]
port 207 nsew signal bidirectional
rlabel metal3 s 0 55028 800 55268 6 wbs_dat_o[30]
port 208 nsew signal bidirectional
rlabel metal3 s 69200 50948 70000 51188 6 wbs_dat_o[31]
port 209 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 wbs_dat_o[3]
port 210 nsew signal bidirectional
rlabel metal2 s 24462 0 24574 800 6 wbs_dat_o[4]
port 211 nsew signal bidirectional
rlabel metal2 s 39918 0 40030 800 6 wbs_dat_o[5]
port 212 nsew signal bidirectional
rlabel metal3 s 69200 49588 70000 49828 6 wbs_dat_o[6]
port 213 nsew signal bidirectional
rlabel metal2 s 41206 0 41318 800 6 wbs_dat_o[7]
port 214 nsew signal bidirectional
rlabel metal2 s 48934 71200 49046 72000 6 wbs_dat_o[8]
port 215 nsew signal bidirectional
rlabel metal2 s 47646 71200 47758 72000 6 wbs_dat_o[9]
port 216 nsew signal bidirectional
rlabel metal3 s 0 69988 800 70228 6 wbs_sel_i[0]
port 217 nsew signal input
rlabel metal2 s 10294 71200 10406 72000 6 wbs_sel_i[1]
port 218 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 wbs_sel_i[2]
port 219 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 wbs_sel_i[3]
port 220 nsew signal input
rlabel metal3 s 0 60468 800 60708 6 wbs_stb_i
port 221 nsew signal input
rlabel metal3 s 69200 33948 70000 34188 6 wbs_we_i
port 222 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 72000
<< end >>
