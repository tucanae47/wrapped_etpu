magic
tech sky130A
magscale 1 2
timestamp 1654694708
<< obsli1 >>
rect 1104 2159 68816 69649
<< obsm1 >>
rect 842 2128 68986 69680
<< metal2 >>
rect 634 71200 746 72000
rect 1922 71200 2034 72000
rect 3210 71200 3322 72000
rect 4498 71200 4610 72000
rect 5786 71200 5898 72000
rect 7074 71200 7186 72000
rect 8362 71200 8474 72000
rect 9650 71200 9762 72000
rect 10938 71200 11050 72000
rect 12226 71200 12338 72000
rect 13514 71200 13626 72000
rect 14802 71200 14914 72000
rect 16090 71200 16202 72000
rect 17378 71200 17490 72000
rect 18666 71200 18778 72000
rect 19954 71200 20066 72000
rect 21242 71200 21354 72000
rect 22530 71200 22642 72000
rect 24462 71200 24574 72000
rect 25750 71200 25862 72000
rect 27038 71200 27150 72000
rect 28326 71200 28438 72000
rect 29614 71200 29726 72000
rect 30902 71200 31014 72000
rect 32190 71200 32302 72000
rect 33478 71200 33590 72000
rect 34766 71200 34878 72000
rect 36054 71200 36166 72000
rect 37342 71200 37454 72000
rect 38630 71200 38742 72000
rect 39918 71200 40030 72000
rect 41206 71200 41318 72000
rect 42494 71200 42606 72000
rect 43782 71200 43894 72000
rect 45070 71200 45182 72000
rect 46358 71200 46470 72000
rect 47646 71200 47758 72000
rect 48934 71200 49046 72000
rect 50222 71200 50334 72000
rect 51510 71200 51622 72000
rect 52798 71200 52910 72000
rect 54086 71200 54198 72000
rect 55374 71200 55486 72000
rect 56662 71200 56774 72000
rect 57950 71200 58062 72000
rect 59238 71200 59350 72000
rect 60526 71200 60638 72000
rect 61814 71200 61926 72000
rect 63102 71200 63214 72000
rect 64390 71200 64502 72000
rect 65678 71200 65790 72000
rect 66966 71200 67078 72000
rect 68254 71200 68366 72000
rect 69542 71200 69654 72000
rect -10 0 102 800
rect 1278 0 1390 800
rect 2566 0 2678 800
rect 3854 0 3966 800
rect 5142 0 5254 800
rect 6430 0 6542 800
rect 7718 0 7830 800
rect 9006 0 9118 800
rect 10294 0 10406 800
rect 11582 0 11694 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 15446 0 15558 800
rect 16734 0 16846 800
rect 18022 0 18134 800
rect 19310 0 19422 800
rect 20598 0 20710 800
rect 21886 0 21998 800
rect 23174 0 23286 800
rect 24462 0 24574 800
rect 25750 0 25862 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 29614 0 29726 800
rect 30902 0 31014 800
rect 32190 0 32302 800
rect 33478 0 33590 800
rect 34766 0 34878 800
rect 36054 0 36166 800
rect 37342 0 37454 800
rect 38630 0 38742 800
rect 39918 0 40030 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43782 0 43894 800
rect 45070 0 45182 800
rect 47002 0 47114 800
rect 48290 0 48402 800
rect 49578 0 49690 800
rect 50866 0 50978 800
rect 52154 0 52266 800
rect 53442 0 53554 800
rect 54730 0 54842 800
rect 56018 0 56130 800
rect 57306 0 57418 800
rect 58594 0 58706 800
rect 59882 0 59994 800
rect 61170 0 61282 800
rect 62458 0 62570 800
rect 63746 0 63858 800
rect 65034 0 65146 800
rect 66322 0 66434 800
rect 67610 0 67722 800
rect 68898 0 69010 800
<< obsm2 >>
rect 848 71144 1866 71346
rect 2090 71144 3154 71346
rect 3378 71144 4442 71346
rect 4666 71144 5730 71346
rect 5954 71144 7018 71346
rect 7242 71144 8306 71346
rect 8530 71144 9594 71346
rect 9818 71144 10882 71346
rect 11106 71144 12170 71346
rect 12394 71144 13458 71346
rect 13682 71144 14746 71346
rect 14970 71144 16034 71346
rect 16258 71144 17322 71346
rect 17546 71144 18610 71346
rect 18834 71144 19898 71346
rect 20122 71144 21186 71346
rect 21410 71144 22474 71346
rect 22698 71144 24406 71346
rect 24630 71144 25694 71346
rect 25918 71144 26982 71346
rect 27206 71144 28270 71346
rect 28494 71144 29558 71346
rect 29782 71144 30846 71346
rect 31070 71144 32134 71346
rect 32358 71144 33422 71346
rect 33646 71144 34710 71346
rect 34934 71144 35998 71346
rect 36222 71144 37286 71346
rect 37510 71144 38574 71346
rect 38798 71144 39862 71346
rect 40086 71144 41150 71346
rect 41374 71144 42438 71346
rect 42662 71144 43726 71346
rect 43950 71144 45014 71346
rect 45238 71144 46302 71346
rect 46526 71144 47590 71346
rect 47814 71144 48878 71346
rect 49102 71144 50166 71346
rect 50390 71144 51454 71346
rect 51678 71144 52742 71346
rect 52966 71144 54030 71346
rect 54254 71144 55318 71346
rect 55542 71144 56606 71346
rect 56830 71144 57894 71346
rect 58118 71144 59182 71346
rect 59406 71144 60470 71346
rect 60694 71144 61758 71346
rect 61982 71144 63046 71346
rect 63270 71144 64334 71346
rect 64558 71144 65622 71346
rect 65846 71144 66910 71346
rect 67134 71144 68198 71346
rect 68422 71144 68980 71346
rect 848 856 68980 71144
rect 848 734 1222 856
rect 1446 734 2510 856
rect 2734 734 3798 856
rect 4022 734 5086 856
rect 5310 734 6374 856
rect 6598 734 7662 856
rect 7886 734 8950 856
rect 9174 734 10238 856
rect 10462 734 11526 856
rect 11750 734 12814 856
rect 13038 734 14102 856
rect 14326 734 15390 856
rect 15614 734 16678 856
rect 16902 734 17966 856
rect 18190 734 19254 856
rect 19478 734 20542 856
rect 20766 734 21830 856
rect 22054 734 23118 856
rect 23342 734 24406 856
rect 24630 734 25694 856
rect 25918 734 26982 856
rect 27206 734 28270 856
rect 28494 734 29558 856
rect 29782 734 30846 856
rect 31070 734 32134 856
rect 32358 734 33422 856
rect 33646 734 34710 856
rect 34934 734 35998 856
rect 36222 734 37286 856
rect 37510 734 38574 856
rect 38798 734 39862 856
rect 40086 734 41150 856
rect 41374 734 42438 856
rect 42662 734 43726 856
rect 43950 734 45014 856
rect 45238 734 46946 856
rect 47170 734 48234 856
rect 48458 734 49522 856
rect 49746 734 50810 856
rect 51034 734 52098 856
rect 52322 734 53386 856
rect 53610 734 54674 856
rect 54898 734 55962 856
rect 56186 734 57250 856
rect 57474 734 58538 856
rect 58762 734 59826 856
rect 60050 734 61114 856
rect 61338 734 62402 856
rect 62626 734 63690 856
rect 63914 734 64978 856
rect 65202 734 66266 856
rect 66490 734 67554 856
rect 67778 734 68842 856
<< metal3 >>
rect 0 71348 800 71588
rect 0 69988 800 70228
rect 69200 69988 70000 70228
rect 0 68628 800 68868
rect 69200 68628 70000 68868
rect 0 67268 800 67508
rect 69200 67268 70000 67508
rect 0 65908 800 66148
rect 69200 65908 70000 66148
rect 0 64548 800 64788
rect 69200 64548 70000 64788
rect 0 63188 800 63428
rect 69200 63188 70000 63428
rect 0 61828 800 62068
rect 69200 61828 70000 62068
rect 0 60468 800 60708
rect 69200 60468 70000 60708
rect 0 59108 800 59348
rect 69200 59108 70000 59348
rect 0 57748 800 57988
rect 69200 57748 70000 57988
rect 0 56388 800 56628
rect 69200 56388 70000 56628
rect 0 55028 800 55268
rect 69200 55028 70000 55268
rect 0 53668 800 53908
rect 69200 53668 70000 53908
rect 0 52308 800 52548
rect 69200 52308 70000 52548
rect 0 50948 800 51188
rect 69200 50948 70000 51188
rect 0 49588 800 49828
rect 69200 49588 70000 49828
rect 69200 48228 70000 48468
rect 0 47548 800 47788
rect 69200 46868 70000 47108
rect 0 46188 800 46428
rect 69200 45508 70000 45748
rect 0 44828 800 45068
rect 69200 44148 70000 44388
rect 0 43468 800 43708
rect 69200 42788 70000 43028
rect 0 42108 800 42348
rect 69200 41428 70000 41668
rect 0 40748 800 40988
rect 69200 40068 70000 40308
rect 0 39388 800 39628
rect 69200 38708 70000 38948
rect 0 38028 800 38268
rect 69200 37348 70000 37588
rect 0 36668 800 36908
rect 69200 35988 70000 36228
rect 0 35308 800 35548
rect 69200 34628 70000 34868
rect 0 33948 800 34188
rect 69200 33268 70000 33508
rect 0 32588 800 32828
rect 69200 31908 70000 32148
rect 0 31228 800 31468
rect 69200 30548 70000 30788
rect 0 29868 800 30108
rect 69200 29188 70000 29428
rect 0 28508 800 28748
rect 69200 27828 70000 28068
rect 0 27148 800 27388
rect 69200 26468 70000 26708
rect 0 25788 800 26028
rect 69200 25108 70000 25348
rect 0 24428 800 24668
rect 69200 23748 70000 23988
rect 0 23068 800 23308
rect 0 21708 800 21948
rect 69200 21708 70000 21948
rect 0 20348 800 20588
rect 69200 20348 70000 20588
rect 0 18988 800 19228
rect 69200 18988 70000 19228
rect 0 17628 800 17868
rect 69200 17628 70000 17868
rect 0 16268 800 16508
rect 69200 16268 70000 16508
rect 0 14908 800 15148
rect 69200 14908 70000 15148
rect 0 13548 800 13788
rect 69200 13548 70000 13788
rect 0 12188 800 12428
rect 69200 12188 70000 12428
rect 0 10828 800 11068
rect 69200 10828 70000 11068
rect 0 9468 800 9708
rect 69200 9468 70000 9708
rect 0 8108 800 8348
rect 69200 8108 70000 8348
rect 0 6748 800 6988
rect 69200 6748 70000 6988
rect 0 5388 800 5628
rect 69200 5388 70000 5628
rect 0 4028 800 4268
rect 69200 4028 70000 4268
rect 0 2668 800 2908
rect 69200 2668 70000 2908
rect 0 1308 800 1548
rect 69200 1308 70000 1548
rect 69200 -52 70000 188
<< obsm3 >>
rect 880 69908 69120 70141
rect 800 68948 69200 69908
rect 880 68548 69120 68948
rect 800 67588 69200 68548
rect 880 67188 69120 67588
rect 800 66228 69200 67188
rect 880 65828 69120 66228
rect 800 64868 69200 65828
rect 880 64468 69120 64868
rect 800 63508 69200 64468
rect 880 63108 69120 63508
rect 800 62148 69200 63108
rect 880 61748 69120 62148
rect 800 60788 69200 61748
rect 880 60388 69120 60788
rect 800 59428 69200 60388
rect 880 59028 69120 59428
rect 800 58068 69200 59028
rect 880 57668 69120 58068
rect 800 56708 69200 57668
rect 880 56308 69120 56708
rect 800 55348 69200 56308
rect 880 54948 69120 55348
rect 800 53988 69200 54948
rect 880 53588 69120 53988
rect 800 52628 69200 53588
rect 880 52228 69120 52628
rect 800 51268 69200 52228
rect 880 50868 69120 51268
rect 800 49908 69200 50868
rect 880 49508 69120 49908
rect 800 48548 69200 49508
rect 800 48148 69120 48548
rect 800 47868 69200 48148
rect 880 47468 69200 47868
rect 800 47188 69200 47468
rect 800 46788 69120 47188
rect 800 46508 69200 46788
rect 880 46108 69200 46508
rect 800 45828 69200 46108
rect 800 45428 69120 45828
rect 800 45148 69200 45428
rect 880 44748 69200 45148
rect 800 44468 69200 44748
rect 800 44068 69120 44468
rect 800 43788 69200 44068
rect 880 43388 69200 43788
rect 800 43108 69200 43388
rect 800 42708 69120 43108
rect 800 42428 69200 42708
rect 880 42028 69200 42428
rect 800 41748 69200 42028
rect 800 41348 69120 41748
rect 800 41068 69200 41348
rect 880 40668 69200 41068
rect 800 40388 69200 40668
rect 800 39988 69120 40388
rect 800 39708 69200 39988
rect 880 39308 69200 39708
rect 800 39028 69200 39308
rect 800 38628 69120 39028
rect 800 38348 69200 38628
rect 880 37948 69200 38348
rect 800 37668 69200 37948
rect 800 37268 69120 37668
rect 800 36988 69200 37268
rect 880 36588 69200 36988
rect 800 36308 69200 36588
rect 800 35908 69120 36308
rect 800 35628 69200 35908
rect 880 35228 69200 35628
rect 800 34948 69200 35228
rect 800 34548 69120 34948
rect 800 34268 69200 34548
rect 880 33868 69200 34268
rect 800 33588 69200 33868
rect 800 33188 69120 33588
rect 800 32908 69200 33188
rect 880 32508 69200 32908
rect 800 32228 69200 32508
rect 800 31828 69120 32228
rect 800 31548 69200 31828
rect 880 31148 69200 31548
rect 800 30868 69200 31148
rect 800 30468 69120 30868
rect 800 30188 69200 30468
rect 880 29788 69200 30188
rect 800 29508 69200 29788
rect 800 29108 69120 29508
rect 800 28828 69200 29108
rect 880 28428 69200 28828
rect 800 28148 69200 28428
rect 800 27748 69120 28148
rect 800 27468 69200 27748
rect 880 27068 69200 27468
rect 800 26788 69200 27068
rect 800 26388 69120 26788
rect 800 26108 69200 26388
rect 880 25708 69200 26108
rect 800 25428 69200 25708
rect 800 25028 69120 25428
rect 800 24748 69200 25028
rect 880 24348 69200 24748
rect 800 24068 69200 24348
rect 800 23668 69120 24068
rect 800 23388 69200 23668
rect 880 22988 69200 23388
rect 800 22028 69200 22988
rect 880 21628 69120 22028
rect 800 20668 69200 21628
rect 880 20268 69120 20668
rect 800 19308 69200 20268
rect 880 18908 69120 19308
rect 800 17948 69200 18908
rect 880 17548 69120 17948
rect 800 16588 69200 17548
rect 880 16188 69120 16588
rect 800 15228 69200 16188
rect 880 14828 69120 15228
rect 800 13868 69200 14828
rect 880 13468 69120 13868
rect 800 12508 69200 13468
rect 880 12108 69120 12508
rect 800 11148 69200 12108
rect 880 10748 69120 11148
rect 800 9788 69200 10748
rect 880 9388 69120 9788
rect 800 8428 69200 9388
rect 880 8028 69120 8428
rect 800 7068 69200 8028
rect 880 6668 69120 7068
rect 800 5708 69200 6668
rect 880 5308 69120 5708
rect 800 4348 69200 5308
rect 880 3948 69120 4348
rect 800 2988 69200 3948
rect 880 2588 69120 2988
rect 800 1628 69200 2588
rect 880 1395 69120 1628
<< metal4 >>
rect 4208 2128 4528 69680
rect 19568 2128 19888 69680
rect 34928 2128 35248 69680
rect 50288 2128 50608 69680
rect 65648 2128 65968 69680
<< labels >>
rlabel metal3 s 0 65908 800 66148 6 active
port 1 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 38630 71200 38742 72000 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 0 71348 800 71588 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 69200 60468 70000 60708 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 33478 0 33590 800 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 25750 71200 25862 72000 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 69200 63188 70000 63428 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 69200 6748 70000 6988 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 13514 71200 13626 72000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 16090 71200 16202 72000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 61170 0 61282 800 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 69200 23748 70000 23988 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 12226 71200 12338 72000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 8362 71200 8474 72000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 53442 0 53554 800 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 52154 0 52266 800 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 69200 16268 70000 16508 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 69542 71200 69654 72000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 69200 29188 70000 29428 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 0 63188 800 63428 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 0 36668 800 36908 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 52798 71200 52910 72000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 60526 71200 60638 72000 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 69200 45508 70000 45748 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 61814 71200 61926 72000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 39918 71200 40030 72000 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 69200 44148 70000 44388 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 69200 68628 70000 68868 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 0 43468 800 43708 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 69200 48228 70000 48468 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 10938 71200 11050 72000 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 io_oeb[0]
port 40 nsew signal bidirectional
rlabel metal3 s 0 24428 800 24668 6 io_oeb[10]
port 41 nsew signal bidirectional
rlabel metal3 s 69200 41428 70000 41668 6 io_oeb[11]
port 42 nsew signal bidirectional
rlabel metal3 s 69200 21708 70000 21948 6 io_oeb[12]
port 43 nsew signal bidirectional
rlabel metal3 s 69200 20348 70000 20588 6 io_oeb[13]
port 44 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 io_oeb[14]
port 45 nsew signal bidirectional
rlabel metal2 s 18666 71200 18778 72000 6 io_oeb[15]
port 46 nsew signal bidirectional
rlabel metal3 s 69200 4028 70000 4268 6 io_oeb[16]
port 47 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 io_oeb[17]
port 48 nsew signal bidirectional
rlabel metal2 s 50222 71200 50334 72000 6 io_oeb[18]
port 49 nsew signal bidirectional
rlabel metal2 s 19954 71200 20066 72000 6 io_oeb[19]
port 50 nsew signal bidirectional
rlabel metal2 s 56018 0 56130 800 6 io_oeb[1]
port 51 nsew signal bidirectional
rlabel metal3 s 69200 31908 70000 32148 6 io_oeb[20]
port 52 nsew signal bidirectional
rlabel metal2 s 1922 71200 2034 72000 6 io_oeb[21]
port 53 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 io_oeb[22]
port 54 nsew signal bidirectional
rlabel metal2 s 34766 71200 34878 72000 6 io_oeb[23]
port 55 nsew signal bidirectional
rlabel metal2 s 36054 71200 36166 72000 6 io_oeb[24]
port 56 nsew signal bidirectional
rlabel metal2 s 67610 0 67722 800 6 io_oeb[25]
port 57 nsew signal bidirectional
rlabel metal3 s 69200 56388 70000 56628 6 io_oeb[26]
port 58 nsew signal bidirectional
rlabel metal2 s 41206 71200 41318 72000 6 io_oeb[27]
port 59 nsew signal bidirectional
rlabel metal2 s 59882 0 59994 800 6 io_oeb[28]
port 60 nsew signal bidirectional
rlabel metal3 s 69200 46868 70000 47108 6 io_oeb[29]
port 61 nsew signal bidirectional
rlabel metal2 s 57950 71200 58062 72000 6 io_oeb[2]
port 62 nsew signal bidirectional
rlabel metal2 s 3210 71200 3322 72000 6 io_oeb[30]
port 63 nsew signal bidirectional
rlabel metal2 s 58594 0 58706 800 6 io_oeb[31]
port 64 nsew signal bidirectional
rlabel metal3 s 0 35308 800 35548 6 io_oeb[32]
port 65 nsew signal bidirectional
rlabel metal2 s 68898 0 69010 800 6 io_oeb[33]
port 66 nsew signal bidirectional
rlabel metal2 s 14802 71200 14914 72000 6 io_oeb[34]
port 67 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 io_oeb[35]
port 68 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 io_oeb[36]
port 69 nsew signal bidirectional
rlabel metal3 s 0 25788 800 26028 6 io_oeb[37]
port 70 nsew signal bidirectional
rlabel metal2 s 36054 0 36166 800 6 io_oeb[3]
port 71 nsew signal bidirectional
rlabel metal3 s 69200 1308 70000 1548 6 io_oeb[4]
port 72 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 io_oeb[5]
port 73 nsew signal bidirectional
rlabel metal3 s 69200 26468 70000 26708 6 io_oeb[6]
port 74 nsew signal bidirectional
rlabel metal2 s 17378 71200 17490 72000 6 io_oeb[7]
port 75 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 io_oeb[8]
port 76 nsew signal bidirectional
rlabel metal2 s 15446 0 15558 800 6 io_oeb[9]
port 77 nsew signal bidirectional
rlabel metal3 s 69200 67268 70000 67508 6 io_out[0]
port 78 nsew signal bidirectional
rlabel metal3 s 69200 40068 70000 40308 6 io_out[10]
port 79 nsew signal bidirectional
rlabel metal3 s 0 4028 800 4268 6 io_out[11]
port 80 nsew signal bidirectional
rlabel metal3 s 0 10828 800 11068 6 io_out[12]
port 81 nsew signal bidirectional
rlabel metal2 s 57306 0 57418 800 6 io_out[13]
port 82 nsew signal bidirectional
rlabel metal3 s 69200 57748 70000 57988 6 io_out[14]
port 83 nsew signal bidirectional
rlabel metal3 s 0 59108 800 59348 6 io_out[15]
port 84 nsew signal bidirectional
rlabel metal3 s 69200 38708 70000 38948 6 io_out[16]
port 85 nsew signal bidirectional
rlabel metal2 s 64390 71200 64502 72000 6 io_out[17]
port 86 nsew signal bidirectional
rlabel metal2 s 66322 0 66434 800 6 io_out[18]
port 87 nsew signal bidirectional
rlabel metal3 s 0 33948 800 34188 6 io_out[19]
port 88 nsew signal bidirectional
rlabel metal2 s 46358 71200 46470 72000 6 io_out[1]
port 89 nsew signal bidirectional
rlabel metal2 s 56662 71200 56774 72000 6 io_out[20]
port 90 nsew signal bidirectional
rlabel metal3 s 0 57748 800 57988 6 io_out[21]
port 91 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 io_out[22]
port 92 nsew signal bidirectional
rlabel metal3 s 69200 33268 70000 33508 6 io_out[23]
port 93 nsew signal bidirectional
rlabel metal2 s 38630 0 38742 800 6 io_out[24]
port 94 nsew signal bidirectional
rlabel metal2 s 51510 71200 51622 72000 6 io_out[25]
port 95 nsew signal bidirectional
rlabel metal3 s 0 8108 800 8348 6 io_out[26]
port 96 nsew signal bidirectional
rlabel metal2 s 54086 71200 54198 72000 6 io_out[27]
port 97 nsew signal bidirectional
rlabel metal2 s 24462 0 24574 800 6 io_out[28]
port 98 nsew signal bidirectional
rlabel metal3 s 69200 2668 70000 2908 6 io_out[29]
port 99 nsew signal bidirectional
rlabel metal2 s 10294 0 10406 800 6 io_out[2]
port 100 nsew signal bidirectional
rlabel metal3 s 0 9468 800 9708 6 io_out[30]
port 101 nsew signal bidirectional
rlabel metal3 s 0 20348 800 20588 6 io_out[31]
port 102 nsew signal bidirectional
rlabel metal3 s 0 67268 800 67508 6 io_out[32]
port 103 nsew signal bidirectional
rlabel metal3 s 69200 10828 70000 11068 6 io_out[33]
port 104 nsew signal bidirectional
rlabel metal3 s 69200 59108 70000 59348 6 io_out[34]
port 105 nsew signal bidirectional
rlabel metal3 s 69200 55028 70000 55268 6 io_out[35]
port 106 nsew signal bidirectional
rlabel metal2 s 21242 71200 21354 72000 6 io_out[36]
port 107 nsew signal bidirectional
rlabel metal3 s 69200 64548 70000 64788 6 io_out[37]
port 108 nsew signal bidirectional
rlabel metal3 s 0 61828 800 62068 6 io_out[3]
port 109 nsew signal bidirectional
rlabel metal3 s 69200 42788 70000 43028 6 io_out[4]
port 110 nsew signal bidirectional
rlabel metal2 s 32190 71200 32302 72000 6 io_out[5]
port 111 nsew signal bidirectional
rlabel metal2 s 66966 71200 67078 72000 6 io_out[6]
port 112 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 io_out[7]
port 113 nsew signal bidirectional
rlabel metal2 s 27038 0 27150 800 6 io_out[8]
port 114 nsew signal bidirectional
rlabel metal3 s 0 21708 800 21948 6 io_out[9]
port 115 nsew signal bidirectional
rlabel metal3 s 69200 12188 70000 12428 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 30902 0 31014 800 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 69200 9468 70000 9708 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 53668 800 53908 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 18988 800 19228 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal2 s 22530 71200 22642 72000 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 43782 71200 43894 72000 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal2 s 33478 71200 33590 72000 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal2 s 62458 0 62570 800 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 24462 71200 24574 72000 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 52308 800 52548 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal2 s 68254 71200 68366 72000 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 69200 13548 70000 13788 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 1308 800 1548 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 55028 800 55268 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 69200 5388 70000 5628 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal2 s 634 71200 746 72000 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal2 s 54730 0 54842 800 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 59238 71200 59350 72000 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 69200 35988 70000 36228 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 27038 71200 27150 72000 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 28326 71200 28438 72000 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_data_out[0]
port 148 nsew signal bidirectional
rlabel metal3 s 69200 17628 70000 17868 6 la1_data_out[10]
port 149 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la1_data_out[11]
port 150 nsew signal bidirectional
rlabel metal3 s 69200 65908 70000 66148 6 la1_data_out[12]
port 151 nsew signal bidirectional
rlabel metal2 s 5786 71200 5898 72000 6 la1_data_out[13]
port 152 nsew signal bidirectional
rlabel metal2 s 37342 71200 37454 72000 6 la1_data_out[14]
port 153 nsew signal bidirectional
rlabel metal3 s 0 2668 800 2908 6 la1_data_out[15]
port 154 nsew signal bidirectional
rlabel metal3 s 69200 25108 70000 25348 6 la1_data_out[16]
port 155 nsew signal bidirectional
rlabel metal3 s 69200 52308 70000 52548 6 la1_data_out[17]
port 156 nsew signal bidirectional
rlabel metal2 s 7074 71200 7186 72000 6 la1_data_out[18]
port 157 nsew signal bidirectional
rlabel metal3 s 69200 37348 70000 37588 6 la1_data_out[19]
port 158 nsew signal bidirectional
rlabel metal3 s 0 64548 800 64788 6 la1_data_out[1]
port 159 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la1_data_out[20]
port 160 nsew signal bidirectional
rlabel metal3 s 69200 61828 70000 62068 6 la1_data_out[21]
port 161 nsew signal bidirectional
rlabel metal2 s 42494 71200 42606 72000 6 la1_data_out[22]
port 162 nsew signal bidirectional
rlabel metal2 s 18022 0 18134 800 6 la1_data_out[23]
port 163 nsew signal bidirectional
rlabel metal3 s 69200 27828 70000 28068 6 la1_data_out[24]
port 164 nsew signal bidirectional
rlabel metal3 s 0 5388 800 5628 6 la1_data_out[25]
port 165 nsew signal bidirectional
rlabel metal3 s 69200 8108 70000 8348 6 la1_data_out[26]
port 166 nsew signal bidirectional
rlabel metal3 s 0 68628 800 68868 6 la1_data_out[27]
port 167 nsew signal bidirectional
rlabel metal2 s 63746 0 63858 800 6 la1_data_out[28]
port 168 nsew signal bidirectional
rlabel metal2 s 9006 0 9118 800 6 la1_data_out[29]
port 169 nsew signal bidirectional
rlabel metal2 s 29614 0 29726 800 6 la1_data_out[2]
port 170 nsew signal bidirectional
rlabel metal3 s 69200 18988 70000 19228 6 la1_data_out[30]
port 171 nsew signal bidirectional
rlabel metal3 s 69200 69988 70000 70228 6 la1_data_out[31]
port 172 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la1_data_out[3]
port 173 nsew signal bidirectional
rlabel metal2 s 65034 0 65146 800 6 la1_data_out[4]
port 174 nsew signal bidirectional
rlabel metal2 s 5142 0 5254 800 6 la1_data_out[5]
port 175 nsew signal bidirectional
rlabel metal3 s 69200 30548 70000 30788 6 la1_data_out[6]
port 176 nsew signal bidirectional
rlabel metal2 s 1278 0 1390 800 6 la1_data_out[7]
port 177 nsew signal bidirectional
rlabel metal3 s 69200 53668 70000 53908 6 la1_data_out[8]
port 178 nsew signal bidirectional
rlabel metal2 s 65678 71200 65790 72000 6 la1_data_out[9]
port 179 nsew signal bidirectional
rlabel metal3 s 69200 -52 70000 188 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal2 s 63102 71200 63214 72000 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal2 s 42494 0 42606 800 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 50866 0 50978 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 0 50948 800 51188 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal2 s 4498 71200 4610 72000 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 30902 71200 31014 72000 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal2 s 3854 0 3966 800 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal2 s 45070 71200 45182 72000 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 29614 71200 29726 72000 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal2 s 55374 71200 55486 72000 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 69200 14908 70000 15148 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 0 56388 800 56628 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 69200 50948 70000 51188 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 69200 49588 70000 49828 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 48934 71200 49046 72000 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal2 s 47646 71200 47758 72000 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 0 69988 800 70228 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal2 s 9650 71200 9762 72000 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 0 60468 800 60708 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 2128 4528 69680 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 2128 35248 69680 6 vccd1
port 212 nsew power input
rlabel metal4 s 65648 2128 65968 69680 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 2128 19888 69680 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 2128 50608 69680 6 vssd1
port 213 nsew ground input
rlabel metal3 s 69200 34628 70000 34868 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 72000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1802336
string GDS_FILE /home/tuc/MPW5/caravel_user_project/openlane/wrapped_etpu/runs/wrapped_etpu/results/finishing/wrapped_etpu.magic.gds
string GDS_START 77506
<< end >>

